// [5:0]AxUSER driven by PL-AXI_ID
// [15:6]AxUSER need to be tied to 10'b0000001111

module RawPS8(

// ps_to_pl supplied by PS to the PL
// pl_to_ps supplied by PL to the PS

// Clocks (all unbuffered)
output wire clk_ps_to_pl_dp_video,
output wire clk_ps_to_pl_dp_audio,
output wire clk_ps_to_pl_fmio_gem0_fifo_tx,
output wire clk_ps_to_pl_fmio_gem0_fifo_rx,
output wire clk_ps_to_pl_fmio_gem1_fifo_tx,
output wire clk_ps_to_pl_fmio_gem1_fifo_rx,
output wire clk_ps_to_pl_fmio_gem2_fifo_tx,
output wire clk_ps_to_pl_fmio_gem2_fifo_rx,
output wire clk_ps_to_pl_fmio_gem3_fifo_tx,
output wire clk_ps_to_pl_fmio_gem3_fifo_rx,
output wire clk_ps_to_pl_gem_tsu_clk,
output wire clk_ps_to_pl_emio_sdio0,
output wire clk_ps_to_pl_emio_sdio1,
output wire clk_ps_to_pl_trace,
output wire [3:0] clk_ps_to_pl_clks,

// to ps from pl (tps_fpl)
input  wire clk_ps_to_pl_axi_hpm0_fpd, // PS supplier gp0
input  wire clk_ps_to_pl_axi_hpm0_lpd, // PS supplier gp2
input  wire clk_ps_to_pl_axi_hpm1_fpd, // PS supplier gp1
input  wire clk_pl_to_ps_axi_hpc0_fpd_read,  // PS consumer gp0 read
input  wire clk_pl_to_ps_axi_hpc0_fpd_write, // PS consumer gp0 write
input  wire clk_pl_to_ps_axi_hpc1_fpd_read,  // PS consumer gp1 read
input  wire clk_pl_to_ps_axi_hpc1_fpd_write, // PS consumer gp1 write
input  wire clk_pl_to_ps_axi_hp0_fpd_read,   // PS consumer gp2 read
input  wire clk_pl_to_ps_axi_hp0_fpd_write,  // PS consumer gp2 write
input  wire clk_pl_to_ps_axi_hp1_fpd_read,   // PS consumer gp3 read
input  wire clk_pl_to_ps_axi_hp1_fpd_write,  // PS consumer gp3 write
input  wire clk_pl_to_ps_axi_hp2_fpd_read,   // PS consumer gp4 read
input  wire clk_pl_to_ps_axi_hp2_fpd_write,  // PS consumer gp4 write
input  wire clk_pl_to_ps_axi_hp3_fpd_read,   // PS consumer gp5 read
input  wire clk_pl_to_ps_axi_hp3_fpd_write,  // PS consumer gp5 write
input  wire clk_pl_to_ps_axi_lpd_read,       // PS consumer gp6 read
input  wire clk_pl_to_ps_axi_lpd_write,      // PS consumer gp6 write
input  wire clk_pl_to_ps_axi_acp_fpd,        // PS consumer acp
input  wire clk_pl_to_ps_axi_ace_fpd,        // PS consumer ace

input  wire clk_pl_to_ps_emio_enet0_gmii_rx,
input  wire clk_pl_to_ps_emio_enet0_gmii_tx,
input  wire clk_pl_to_ps_emio_enet1_gmii_rx,
input  wire clk_pl_to_ps_emio_enet1_gmii_tx,
input  wire clk_pl_to_ps_emio_enet2_gmii_rx,
input  wire clk_pl_to_ps_emio_enet2_gmii_tx,
input  wire clk_pl_to_ps_emio_enet3_gmii_rx,
input  wire clk_pl_to_ps_emio_enet3_gmii_tx,
input wire  clk_pl_to_ps_fmio_gem0_fifo_tx,
input wire  clk_pl_to_ps_fmio_gem0_fifo_rx,
input wire  clk_pl_to_ps_fmio_gem1_fifo_tx,
input wire  clk_pl_to_ps_fmio_gem1_fifo_rx,
input wire  clk_pl_to_ps_fmio_gem2_fifo_tx,
input wire  clk_pl_to_ps_fmio_gem2_fifo_rx,
input wire  clk_pl_to_ps_fmio_gem3_fifo_tx,
input wire  clk_pl_to_ps_fmio_gem3_fifo_rx,
input wire  clk_pl_to_ps_fmio_gem_tsu,
input  wire clk_pl_to_ps_emio_enet_tsu,
input  wire clk_pl_to_ps_emio_sdio0,
input  wire clk_pl_to_ps_emio_sdio1,
input wire clk_pl_to_ps_trace,
input  wire [2:0] clk_pl_to_ps_emio_ttc0,
input  wire [2:0] clk_pl_to_ps_emio_ttc1,
input  wire [2:0] clk_pl_to_ps_emio_ttc2,
input  wire [2:0] clk_pl_to_ps_emio_ttc3,
input  wire clk_pl_to_ps_emio_wdt0,
input  wire clk_pl_to_ps_emio_wdt1,
input  wire [7:0] clk_pl_to_ps_adma_fci,
input  wire [7:0] clk_pl_to_ps_gdma_perif,
input  wire [1:0] clk_pl_to_ps_pll_aux_lpd,
input  wire [2:0] clk_pl_to_ps_pll_aux_fpd,
input  wire clk_pl_to_ps_dp_s_axis_audio,
input  wire clk_pl_to_ps_dp_video_in,
input  wire clk_pl_to_ps_ddrc_refresh,
input  [3:0]  clk_pl_to_ps_pstp,

// axi interfaces ports
// 3 128 bit ps to pl axi interfaces
// 8 128 bit pl to ps axi interfaces
output wire [15:0]   ps_to_pl_axi_hpm0_fpd_awid,
output wire [39:0]   ps_to_pl_axi_hpm0_fpd_awaddr,
output wire [7:0]    ps_to_pl_axi_hpm0_fpd_awlen,
output wire [2:0]    ps_to_pl_axi_hpm0_fpd_awsize,
output wire [1:0]    ps_to_pl_axi_hpm0_fpd_awburst,
output wire          ps_to_pl_axi_hpm0_fpd_awlock,
output wire [3:0]    ps_to_pl_axi_hpm0_fpd_awcache,
output wire [2:0]    ps_to_pl_axi_hpm0_fpd_awprot,
output wire          ps_to_pl_axi_hpm0_fpd_awvalid,
output wire [15:0]   ps_to_pl_axi_hpm0_fpd_awuser,
input  wire          ps_to_pl_axi_hpm0_fpd_awready,
output wire [127:0]  ps_to_pl_axi_hpm0_fpd_wdata,
output wire [15:0]   ps_to_pl_axi_hpm0_fpd_wstrb,
output wire          ps_to_pl_axi_hpm0_fpd_wlast,
output wire          ps_to_pl_axi_hpm0_fpd_wvalid,
input  wire          ps_to_pl_axi_hpm0_fpd_wready,
input  wire [15:0]   ps_to_pl_axi_hpm0_fpd_bid,
input  wire [1:0]    ps_to_pl_axi_hpm0_fpd_bresp,
input  wire          ps_to_pl_axi_hpm0_fpd_bvalid,
output wire          ps_to_pl_axi_hpm0_fpd_bready,
output wire [15:0]   ps_to_pl_axi_hpm0_fpd_arid,
output wire [39:0]   ps_to_pl_axi_hpm0_fpd_araddr,
output wire [7:0]    ps_to_pl_axi_hpm0_fpd_arlen,
output wire [2:0]    ps_to_pl_axi_hpm0_fpd_arsize,
output wire [1:0]    ps_to_pl_axi_hpm0_fpd_arburst,
output wire          ps_to_pl_axi_hpm0_fpd_arlock,
output wire [3:0]    ps_to_pl_axi_hpm0_fpd_arcache,
output wire [2:0]    ps_to_pl_axi_hpm0_fpd_arprot,
output wire          ps_to_pl_axi_hpm0_fpd_arvalid,
output wire [15:0]   ps_to_pl_axi_hpm0_fpd_aruser,
input  wire          ps_to_pl_axi_hpm0_fpd_arready,
input  wire [15:0]   ps_to_pl_axi_hpm0_fpd_rid,
input  wire [127:0]  ps_to_pl_axi_hpm0_fpd_rdata,
input  wire [1:0]    ps_to_pl_axi_hpm0_fpd_rresp,
input  wire          ps_to_pl_axi_hpm0_fpd_rlast,
input  wire          ps_to_pl_axi_hpm0_fpd_rvalid,
output wire          ps_to_pl_axi_hpm0_fpd_rready,
output wire [3:0]    ps_to_pl_axi_hpm0_fpd_awqos,
output wire [3:0]    ps_to_pl_axi_hpm0_fpd_arqos,

output wire [15:0]   ps_to_pl_axi_hpm1_fpd_awid,
output wire [39:0]   ps_to_pl_axi_hpm1_fpd_awaddr,
output wire [7:0]    ps_to_pl_axi_hpm1_fpd_awlen,
output wire [2:0]    ps_to_pl_axi_hpm1_fpd_awsize,
output wire [1:0]    ps_to_pl_axi_hpm1_fpd_awburst,
output wire          ps_to_pl_axi_hpm1_fpd_awlock,
output wire [3:0]    ps_to_pl_axi_hpm1_fpd_awcache,
output wire [2:0]    ps_to_pl_axi_hpm1_fpd_awprot,
output wire          ps_to_pl_axi_hpm1_fpd_awvalid,
output wire [15:0]   ps_to_pl_axi_hpm1_fpd_awuser,
input  wire          ps_to_pl_axi_hpm1_fpd_awready,
output wire [127:0]  ps_to_pl_axi_hpm1_fpd_wdata,
output wire [15:0]   ps_to_pl_axi_hpm1_fpd_wstrb,
output wire          ps_to_pl_axi_hpm1_fpd_wlast,
output wire          ps_to_pl_axi_hpm1_fpd_wvalid,
input  wire          ps_to_pl_axi_hpm1_fpd_wready,
input  wire [15:0]   ps_to_pl_axi_hpm1_fpd_bid,
input  wire [1:0]    ps_to_pl_axi_hpm1_fpd_bresp,
input  wire          ps_to_pl_axi_hpm1_fpd_bvalid,
output wire          ps_to_pl_axi_hpm1_fpd_bready,
output wire [15:0]   ps_to_pl_axi_hpm1_fpd_arid,
output wire [39:0]   ps_to_pl_axi_hpm1_fpd_araddr,
output wire [7:0]    ps_to_pl_axi_hpm1_fpd_arlen,
output wire [2:0]    ps_to_pl_axi_hpm1_fpd_arsize,
output wire [1:0]    ps_to_pl_axi_hpm1_fpd_arburst,
output wire          ps_to_pl_axi_hpm1_fpd_arlock,
output wire [3:0]    ps_to_pl_axi_hpm1_fpd_arcache,
output wire [2:0]    ps_to_pl_axi_hpm1_fpd_arprot,
output wire          ps_to_pl_axi_hpm1_fpd_arvalid,
output wire [15:0]   ps_to_pl_axi_hpm1_fpd_aruser,
input  wire          ps_to_pl_axi_hpm1_fpd_arready,
input  wire [15:0]   ps_to_pl_axi_hpm1_fpd_rid,
input  wire [127:0]  ps_to_pl_axi_hpm1_fpd_rdata,
input  wire [1:0]    ps_to_pl_axi_hpm1_fpd_rresp,
input  wire          ps_to_pl_axi_hpm1_fpd_rlast,
input  wire          ps_to_pl_axi_hpm1_fpd_rvalid,
output wire          ps_to_pl_axi_hpm1_fpd_rready,
output wire [3:0]    ps_to_pl_axi_hpm1_fpd_awqos,
output wire [3:0]    ps_to_pl_axi_hpm1_fpd_arqos,

output wire [15:0]   ps_to_pl_axi_hpm0_lpd_awid,
output wire [39:0]   ps_to_pl_axi_hpm0_lpd_awaddr,
output wire [7:0]    ps_to_pl_axi_hpm0_lpd_awlen,
output wire [2:0]    ps_to_pl_axi_hpm0_lpd_awsize,
output wire [1:0]    ps_to_pl_axi_hpm0_lpd_awburst,
output wire          ps_to_pl_axi_hpm0_lpd_awlock,
output wire [3:0]    ps_to_pl_axi_hpm0_lpd_awcache,
output wire [2:0]    ps_to_pl_axi_hpm0_lpd_awprot,
output wire          ps_to_pl_axi_hpm0_lpd_awvalid,
output wire [15:0]   ps_to_pl_axi_hpm0_lpd_awuser,
input  wire          ps_to_pl_axi_hpm0_lpd_awready,
output wire [127:0]  ps_to_pl_axi_hpm0_lpd_wdata,
output wire [15:0]   ps_to_pl_axi_hpm0_lpd_wstrb,
output wire          ps_to_pl_axi_hpm0_lpd_wlast,
output wire          ps_to_pl_axi_hpm0_lpd_wvalid,
input  wire          ps_to_pl_axi_hpm0_lpd_wready,
input  wire [15:0]   ps_to_pl_axi_hpm0_lpd_bid,
input  wire [1:0]    ps_to_pl_axi_hpm0_lpd_bresp,
input  wire          ps_to_pl_axi_hpm0_lpd_bvalid,
output wire          ps_to_pl_axi_hpm0_lpd_bready,
output wire [15:0]   ps_to_pl_axi_hpm0_lpd_arid,
output wire [39:0]   ps_to_pl_axi_hpm0_lpd_araddr,
output wire [7:0]    ps_to_pl_axi_hpm0_lpd_arlen,
output wire [2:0]    ps_to_pl_axi_hpm0_lpd_arsize,
output wire [1:0]    ps_to_pl_axi_hpm0_lpd_arburst,
output wire          ps_to_pl_axi_hpm0_lpd_arlock,
output wire [3:0]    ps_to_pl_axi_hpm0_lpd_arcache,
output wire [2:0]    ps_to_pl_axi_hpm0_lpd_arprot,
output wire          ps_to_pl_axi_hpm0_lpd_arvalid,
output wire [15:0]   ps_to_pl_axi_hpm0_lpd_aruser,
input  wire          ps_to_pl_axi_hpm0_lpd_arready,
input  wire [15:0]   ps_to_pl_axi_hpm0_lpd_rid,
input  wire [127:0]  ps_to_pl_axi_hpm0_lpd_rdata,
input  wire [1:0]    ps_to_pl_axi_hpm0_lpd_rresp,
input  wire          ps_to_pl_axi_hpm0_lpd_rlast,
input  wire          ps_to_pl_axi_hpm0_lpd_rvalid,
output wire          ps_to_pl_axi_hpm0_lpd_rready,
output wire [3:0]    ps_to_pl_axi_hpm0_lpd_awqos,
output wire [3:0]    ps_to_pl_axi_hpm0_lpd_arqos,

input  wire          pl_to_ps_axi_hpc0_fpd_aruser,
input  wire          pl_to_ps_axi_hpc0_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hpc0_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hpc0_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hpc0_fpd_awlen,
input  wire [2:0]    pl_to_ps_axi_hpc0_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hpc0_fpd_awburst,
input  wire          pl_to_ps_axi_hpc0_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hpc0_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hpc0_fpd_awprot,
input  wire          pl_to_ps_axi_hpc0_fpd_awvalid,
output wire          pl_to_ps_axi_hpc0_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hpc0_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hpc0_fpd_wstrb,
input  wire          pl_to_ps_axi_hpc0_fpd_wlast,
input  wire          pl_to_ps_axi_hpc0_fpd_wvalid,
output wire          pl_to_ps_axi_hpc0_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hpc0_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hpc0_fpd_bresp,
output wire          pl_to_ps_axi_hpc0_fpd_bvalid,
input  wire          pl_to_ps_axi_hpc0_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hpc0_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hpc0_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hpc0_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hpc0_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hpc0_fpd_arburst,
input  wire          pl_to_ps_axi_hpc0_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hpc0_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hpc0_fpd_arprot,
input  wire          pl_to_ps_axi_hpc0_fpd_arvalid,
output wire          pl_to_ps_axi_hpc0_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hpc0_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hpc0_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hpc0_fpd_rresp,
output wire          pl_to_ps_axi_hpc0_fpd_rlast,
output wire          pl_to_ps_axi_hpc0_fpd_rvalid,
input  wire          pl_to_ps_axi_hpc0_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hpc0_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hpc0_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hpc0_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hpc0_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hpc0_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hpc0_fpd_wacount,

input  wire          pl_to_ps_axi_hpc1_fpd_aruser,
input  wire          pl_to_ps_axi_hpc1_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hpc1_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hpc1_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hpc1_fpd_awlen,
input  wire [2:0]    pl_to_ps_axi_hpc1_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hpc1_fpd_awburst,
input  wire          pl_to_ps_axi_hpc1_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hpc1_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hpc1_fpd_awprot,
input  wire          pl_to_ps_axi_hpc1_fpd_awvalid,
output wire          pl_to_ps_axi_hpc1_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hpc1_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hpc1_fpd_wstrb,
input  wire          pl_to_ps_axi_hpc1_fpd_wlast,
input  wire          pl_to_ps_axi_hpc1_fpd_wvalid,
output wire          pl_to_ps_axi_hpc1_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hpc1_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hpc1_fpd_bresp,
output wire          pl_to_ps_axi_hpc1_fpd_bvalid,
input  wire          pl_to_ps_axi_hpc1_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hpc1_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hpc1_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hpc1_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hpc1_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hpc1_fpd_arburst,
input  wire          pl_to_ps_axi_hpc1_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hpc1_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hpc1_fpd_arprot,
input  wire          pl_to_ps_axi_hpc1_fpd_arvalid,
output wire          pl_to_ps_axi_hpc1_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hpc1_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hpc1_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hpc1_fpd_rresp,
output wire          pl_to_ps_axi_hpc1_fpd_rlast,
output wire          pl_to_ps_axi_hpc1_fpd_rvalid,
input  wire          pl_to_ps_axi_hpc1_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hpc1_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hpc1_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hpc1_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hpc1_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hpc1_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hpc1_fpd_wacount,

input  wire          pl_to_ps_axi_hp0_fpd_aruser,
input  wire          pl_to_ps_axi_hp0_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hp0_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hp0_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hp0_fpd_awlen ,
input  wire [2:0]    pl_to_ps_axi_hp0_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hp0_fpd_awburst,
input  wire          pl_to_ps_axi_hp0_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hp0_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hp0_fpd_awprot,
input  wire          pl_to_ps_axi_hp0_fpd_awvalid,
output wire          pl_to_ps_axi_hp0_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hp0_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hp0_fpd_wstrb,
input  wire          pl_to_ps_axi_hp0_fpd_wlast,
input  wire          pl_to_ps_axi_hp0_fpd_wvalid,
output wire          pl_to_ps_axi_hp0_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hp0_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hp0_fpd_bresp,
output wire          pl_to_ps_axi_hp0_fpd_bvalid,
input  wire          pl_to_ps_axi_hp0_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hp0_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hp0_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hp0_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hp0_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hp0_fpd_arburst,
input  wire          pl_to_ps_axi_hp0_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hp0_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hp0_fpd_arprot,
input  wire          pl_to_ps_axi_hp0_fpd_arvalid,
output wire          pl_to_ps_axi_hp0_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hp0_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hp0_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hp0_fpd_rresp,
output wire          pl_to_ps_axi_hp0_fpd_rlast,
output wire          pl_to_ps_axi_hp0_fpd_rvalid,
input  wire          pl_to_ps_axi_hp0_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hp0_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hp0_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hp0_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hp0_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hp0_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hp0_fpd_wacount,

input  wire          pl_to_ps_axi_hp1_fpd_aruser,
input  wire          pl_to_ps_axi_hp1_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hp1_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hp1_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hp1_fpd_awlen ,
input  wire [2:0]    pl_to_ps_axi_hp1_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hp1_fpd_awburst,
input  wire          pl_to_ps_axi_hp1_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hp1_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hp1_fpd_awprot,
input  wire          pl_to_ps_axi_hp1_fpd_awvalid,
output wire          pl_to_ps_axi_hp1_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hp1_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hp1_fpd_wstrb,
input  wire          pl_to_ps_axi_hp1_fpd_wlast,
input  wire          pl_to_ps_axi_hp1_fpd_wvalid,
output wire          pl_to_ps_axi_hp1_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hp1_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hp1_fpd_bresp,
output wire          pl_to_ps_axi_hp1_fpd_bvalid,
input  wire          pl_to_ps_axi_hp1_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hp1_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hp1_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hp1_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hp1_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hp1_fpd_arburst,
input  wire          pl_to_ps_axi_hp1_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hp1_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hp1_fpd_arprot,
input  wire          pl_to_ps_axi_hp1_fpd_arvalid,
output wire          pl_to_ps_axi_hp1_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hp1_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hp1_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hp1_fpd_rresp,
output wire          pl_to_ps_axi_hp1_fpd_rlast,
output wire          pl_to_ps_axi_hp1_fpd_rvalid,
input  wire          pl_to_ps_axi_hp1_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hp1_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hp1_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hp1_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hp1_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hp1_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hp1_fpd_wacount,

input  wire          pl_to_ps_axi_hp2_fpd_aruser,
input  wire          pl_to_ps_axi_hp2_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hp2_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hp2_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hp2_fpd_awlen ,
input  wire [2:0]    pl_to_ps_axi_hp2_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hp2_fpd_awburst,
input  wire          pl_to_ps_axi_hp2_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hp2_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hp2_fpd_awprot,
input  wire          pl_to_ps_axi_hp2_fpd_awvalid,
output wire          pl_to_ps_axi_hp2_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hp2_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hp2_fpd_wstrb,
input  wire          pl_to_ps_axi_hp2_fpd_wlast,
input  wire          pl_to_ps_axi_hp2_fpd_wvalid,
output wire          pl_to_ps_axi_hp2_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hp2_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hp2_fpd_bresp,
output wire          pl_to_ps_axi_hp2_fpd_bvalid,
input  wire          pl_to_ps_axi_hp2_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hp2_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hp2_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hp2_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hp2_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hp2_fpd_arburst,
input  wire          pl_to_ps_axi_hp2_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hp2_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hp2_fpd_arprot,
input  wire          pl_to_ps_axi_hp2_fpd_arvalid,
output wire          pl_to_ps_axi_hp2_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hp2_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hp2_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hp2_fpd_rresp,
output wire          pl_to_ps_axi_hp2_fpd_rlast,
output wire          pl_to_ps_axi_hp2_fpd_rvalid,
input  wire          pl_to_ps_axi_hp2_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hp2_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hp2_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hp2_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hp2_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hp2_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hp2_fpd_wacount,

input  wire          pl_to_ps_axi_hp3_fpd_aruser,
input  wire          pl_to_ps_axi_hp3_fpd_awuser,
input  wire [5:0]    pl_to_ps_axi_hp3_fpd_awid,
input  wire [48:0]   pl_to_ps_axi_hp3_fpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_hp3_fpd_awlen ,
input  wire [2:0]    pl_to_ps_axi_hp3_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_hp3_fpd_awburst,
input  wire          pl_to_ps_axi_hp3_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_hp3_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_hp3_fpd_awprot,
input  wire          pl_to_ps_axi_hp3_fpd_awvalid,
output wire          pl_to_ps_axi_hp3_fpd_awready,
input  wire [127:0]  pl_to_ps_axi_hp3_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_hp3_fpd_wstrb,
input  wire          pl_to_ps_axi_hp3_fpd_wlast,
input  wire          pl_to_ps_axi_hp3_fpd_wvalid,
output wire          pl_to_ps_axi_hp3_fpd_wready,
output wire [5:0]    pl_to_ps_axi_hp3_fpd_bid,
output wire [1:0]    pl_to_ps_axi_hp3_fpd_bresp,
output wire          pl_to_ps_axi_hp3_fpd_bvalid,
input  wire          pl_to_ps_axi_hp3_fpd_bready,
input  wire [5:0]    pl_to_ps_axi_hp3_fpd_arid,
input  wire [48:0]   pl_to_ps_axi_hp3_fpd_araddr,
input  wire [7:0]    pl_to_ps_axi_hp3_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_hp3_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_hp3_fpd_arburst,
input  wire          pl_to_ps_axi_hp3_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_hp3_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_hp3_fpd_arprot,
input  wire          pl_to_ps_axi_hp3_fpd_arvalid,
output wire          pl_to_ps_axi_hp3_fpd_arready,
output wire [5:0]    pl_to_ps_axi_hp3_fpd_rid,
output wire [127:0]  pl_to_ps_axi_hp3_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_hp3_fpd_rresp,
output wire          pl_to_ps_axi_hp3_fpd_rlast,
output wire          pl_to_ps_axi_hp3_fpd_rvalid,
input  wire          pl_to_ps_axi_hp3_fpd_rready,
input  wire [3:0]    pl_to_ps_axi_hp3_fpd_awqos,
input  wire [3:0]    pl_to_ps_axi_hp3_fpd_arqos,
output wire [7:0]    pl_to_ps_axi_hp3_fpd_rcount,
output wire [7:0]    pl_to_ps_axi_hp3_fpd_wcount,
output wire [3:0]    pl_to_ps_axi_hp3_fpd_racount,
output wire [3:0]    pl_to_ps_axi_hp3_fpd_wacount,

input  wire          pl_to_ps_axi_lpd_aruser,
input  wire          pl_to_ps_axi_lpd_awuser,
input  wire [5:0]    pl_to_ps_axi_lpd_awid,
input  wire [48:0]   pl_to_ps_axi_lpd_awaddr,
input  wire [7:0]    pl_to_ps_axi_lpd_awlen ,
input  wire [2:0]    pl_to_ps_axi_lpd_awsize,
input  wire [1:0]    pl_to_ps_axi_lpd_awburst,
input  wire          pl_to_ps_axi_lpd_awlock,
input  wire [3:0]    pl_to_ps_axi_lpd_awcache,
input  wire [2:0]    pl_to_ps_axi_lpd_awprot,
input  wire          pl_to_ps_axi_lpd_awvalid,
output wire          pl_to_ps_axi_lpd_awready,
input  wire [127:0]  pl_to_ps_axi_lpd_wdata,
input  wire [15:0]   pl_to_ps_axi_lpd_wstrb,
input  wire          pl_to_ps_axi_lpd_wlast,
input  wire          pl_to_ps_axi_lpd_wvalid,
output wire          pl_to_ps_axi_lpd_wready,
output wire [5:0]    pl_to_ps_axi_lpd_bid,
output wire [1:0]    pl_to_ps_axi_lpd_bresp,
output wire          pl_to_ps_axi_lpd_bvalid,
input  wire          pl_to_ps_axi_lpd_bready,
input  wire [5:0]    pl_to_ps_axi_lpd_arid,
input  wire [48:0]   pl_to_ps_axi_lpd_araddr,
input  wire [7:0]    pl_to_ps_axi_lpd_arlen,
input  wire [2:0]    pl_to_ps_axi_lpd_arsize,
input  wire [1:0]    pl_to_ps_axi_lpd_arburst,
input  wire          pl_to_ps_axi_lpd_arlock,
input  wire [3:0]    pl_to_ps_axi_lpd_arcache,
input  wire [2:0]    pl_to_ps_axi_lpd_arprot,
input  wire          pl_to_ps_axi_lpd_arvalid,
output wire          pl_to_ps_axi_lpd_arready,
output wire [5:0]    pl_to_ps_axi_lpd_rid,
output wire [127:0]  pl_to_ps_axi_lpd_rdata,
output wire [1:0]    pl_to_ps_axi_lpd_rresp,
output wire          pl_to_ps_axi_lpd_rlast,
output wire          pl_to_ps_axi_lpd_rvalid,
input  wire          pl_to_ps_axi_lpd_rready,
input  wire [3:0]    pl_to_ps_axi_lpd_awqos,
input  wire [3:0]    pl_to_ps_axi_lpd_arqos,
output wire [7:0]    pl_to_ps_axi_lpd_rcount,
output wire [7:0]    pl_to_ps_axi_lpd_wcount,
output wire [3:0]    pl_to_ps_axi_lpd_racount,
output wire [3:0]    pl_to_ps_axi_lpd_wacount,

input  wire [39:0]   pl_to_ps_axi_acp_fpd_awaddr,
input  wire [4:0]    pl_to_ps_axi_acp_fpd_awid,
input  wire [7:0]    pl_to_ps_axi_acp_fpd_awlen,
input  wire [2:0]    pl_to_ps_axi_acp_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_acp_fpd_awburst,
input  wire          pl_to_ps_axi_acp_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_acp_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_acp_fpd_awprot,
input  wire          pl_to_ps_axi_acp_fpd_awvalid,
output wire          pl_to_ps_axi_acp_fpd_awready,
input  wire [1:0]    pl_to_ps_axi_acp_fpd_awuser,
input  wire [3:0]    pl_to_ps_axi_acp_fpd_awqos,
input  wire          pl_to_ps_axi_acp_fpd_wlast,
input  wire [127:0]  pl_to_ps_axi_acp_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_acp_fpd_wstrb,
input  wire          pl_to_ps_axi_acp_fpd_wvalid,
output wire          pl_to_ps_axi_acp_fpd_wready,
output wire [1:0]    pl_to_ps_axi_acp_fpd_bresp,
output wire [4:0]    pl_to_ps_axi_acp_fpd_bid,
output wire          pl_to_ps_axi_acp_fpd_bvalid,
input  wire          pl_to_ps_axi_acp_fpd_bready,
input  wire [39:0]   pl_to_ps_axi_acp_fpd_araddr,
input  wire [4:0]    pl_to_ps_axi_acp_fpd_arid,
input  wire [7:0]    pl_to_ps_axi_acp_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_acp_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_acp_fpd_arburst,
input  wire          pl_to_ps_axi_acp_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_acp_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_acp_fpd_arprot,
input  wire          pl_to_ps_axi_acp_fpd_arvalid,
output wire          pl_to_ps_axi_acp_fpd_arready,
input  wire [1:0]    pl_to_ps_axi_acp_fpd_aruser,
input  wire [3:0]    pl_to_ps_axi_acp_fpd_arqos,
output wire [4:0]    pl_to_ps_axi_acp_fpd_rid,
output wire          pl_to_ps_axi_acp_fpd_rlast,
output wire [127:0]  pl_to_ps_axi_acp_fpd_rdata,
output wire [1:0]    pl_to_ps_axi_acp_fpd_rresp,
output wire          pl_to_ps_axi_acp_fpd_rvalid,
input  wire          pl_to_ps_axi_acp_fpd_rready,

input  wire [15:0]   pl_to_ps_axi_ace_fpd_awuser,
input  wire [15:0]   pl_to_ps_axi_ace_fpd_aruser,
input  wire          pl_to_ps_axi_ace_fpd_awvalid,
output wire          pl_to_ps_axi_ace_fpd_awready,
input  wire [5:0]    pl_to_ps_axi_ace_fpd_awid,
input  wire [43:0]   pl_to_ps_axi_ace_fpd_awaddr,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_awregion,
input  wire [7:0]    pl_to_ps_axi_ace_fpd_awlen,
input  wire [2:0]    pl_to_ps_axi_ace_fpd_awsize,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_awburst,
input  wire          pl_to_ps_axi_ace_fpd_awlock,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_awcache,
input  wire [2:0]    pl_to_ps_axi_ace_fpd_awprot,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_awdomain,
input  wire [2:0]    pl_to_ps_axi_ace_fpd_awsnoop,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_awbar,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_awqos,
input  wire          pl_to_ps_axi_ace_fpd_wvalid,
output wire          pl_to_ps_axi_ace_fpd_wready,
input  wire [127:0]  pl_to_ps_axi_ace_fpd_wdata,
input  wire [15:0]   pl_to_ps_axi_ace_fpd_wstrb,
input  wire          pl_to_ps_axi_ace_fpd_wlast,
input  wire          pl_to_ps_axi_ace_fpd_wuser,
output wire          pl_to_ps_axi_ace_fpd_bvalid,
input  wire          pl_to_ps_axi_ace_fpd_bready,
output wire [5:0]    pl_to_ps_axi_ace_fpd_bid,
output wire [1:0]    pl_to_ps_axi_ace_fpd_bresp,
output wire          pl_to_ps_axi_ace_fpd_buser,
input  wire          pl_to_ps_axi_ace_fpd_arvalid,
output wire          pl_to_ps_axi_ace_fpd_arready,
input  wire [5:0]    pl_to_ps_axi_ace_fpd_arid,
input  wire [43:0]   pl_to_ps_axi_ace_fpd_araddr,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_arregion,
input  wire [7:0]    pl_to_ps_axi_ace_fpd_arlen,
input  wire [2:0]    pl_to_ps_axi_ace_fpd_arsize,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_arburst,
input  wire          pl_to_ps_axi_ace_fpd_arlock,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_arcache,
input  wire [2:0]    pl_to_ps_axi_ace_fpd_arprot,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_ardomain,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_arsnoop,
input  wire [1:0]    pl_to_ps_axi_ace_fpd_arbar,
input  wire [3:0]    pl_to_ps_axi_ace_fpd_arqos,
output wire          pl_to_ps_axi_ace_fpd_rvalid,
input  wire          pl_to_ps_axi_ace_fpd_rready,
output wire [5:0]    pl_to_ps_axi_ace_fpd_rid,
output wire [127:0]  pl_to_ps_axi_ace_fpd_rdata,
output wire [3:0]    pl_to_ps_axi_ace_fpd_rresp,
output wire          pl_to_ps_axi_ace_fpd_rlast,
output wire          pl_to_ps_axi_ace_fpd_ruser,
output wire          pl_to_ps_axi_ace_fpd_acvalid,
input  wire          pl_to_ps_axi_ace_fpd_acready,
output wire [43:0]   pl_to_ps_axi_ace_fpd_acaddr,
output wire [3:0]    pl_to_ps_axi_ace_fpd_acsnoop,
output wire [2:0]    pl_to_ps_axi_ace_fpd_acprot,
input  wire          pl_to_ps_axi_ace_fpd_crvalid,
output wire          pl_to_ps_axi_ace_fpd_crready,
input  wire [4:0]    pl_to_ps_axi_ace_fpd_crresp,
input  wire          pl_to_ps_axi_ace_fpd_cdvalid,
output wire          pl_to_ps_axi_ace_fpd_cdready,
input  wire [127:0]  pl_to_ps_axi_ace_fpd_cddata,
input  wire          pl_to_ps_axi_ace_fpd_cdlast,
input  wire          pl_to_ps_axi_ace_fpd_wack,
input  wire          pl_to_ps_axi_ace_fpd_rack,

// supplier and consumer dp audio axi streams
input  wire [31:0] pl_to_ps_axi_stream_dp_audio_tdata,
input  wire pl_to_ps_axi_stream_dp_audio_tid,
input  wire pl_to_ps_axi_stream_dp_audio_tvalid,
output wire pl_to_ps_axi_stream_dp_audio_tready,
output wire [31:0] ps_to_pl_axi_stream_dp_mixed_audio_tdata,
output wire ps_to_pl_axi_stream_dp_mixed_audio_tid,
output wire ps_to_pl_axi_stream_dp_mixed_audio_tvalid,
input  wire ps_to_pl_axi_stream_dp_mixed_audio_tready,


// emio ports
output wire emio_can0_phy_tx,
input  wire emio_can0_phy_rx,

output wire emio_can1_phy_tx,
input  wire emio_can1_phy_rx,

output wire [2:0] emio_enet0_speed_mode,
input  wire emio_enet0_gmii_crs,
input  wire emio_enet0_gmii_col,
input  wire [7:0] emio_enet0_gmii_rxd,
input  wire emio_enet0_gmii_rx_er,
input  wire emio_enet0_gmii_rx_dv,
output wire [7:0] emio_enet0_gmii_txd,
output wire emio_enet0_gmii_tx_en,
output wire emio_enet0_gmii_tx_er,
output wire emio_enet0_mdio_mdc,
input  wire emio_enet0_mdio_i,
output wire emio_enet0_mdio_o,
output wire emio_enet0_mdio_t_n,

output wire [2:0] emio_enet1_speed_mode,
input  wire emio_enet1_gmii_crs,
input  wire emio_enet1_gmii_col,
input  wire [7:0] emio_enet1_gmii_rxd,
input  wire emio_enet1_gmii_rx_er,
input  wire emio_enet1_gmii_rx_dv,
output wire [7:0] emio_enet1_gmii_txd,
output wire emio_enet1_gmii_tx_en,
output wire emio_enet1_gmii_tx_er,
output wire emio_enet1_mdio_mdc,
input  wire emio_enet1_mdio_i,
output wire emio_enet1_mdio_o,
output wire emio_enet1_mdio_t_n,

output wire [2:0] emio_enet2_speed_mode,
input  wire emio_enet2_gmii_crs,
input  wire emio_enet2_gmii_col,
input  wire [7:0] emio_enet2_gmii_rxd,
input  wire emio_enet2_gmii_rx_er,
input  wire emio_enet2_gmii_rx_dv,
output wire [7:0] emio_enet2_gmii_txd,
output wire emio_enet2_gmii_tx_en,
output wire emio_enet2_gmii_tx_er,
output wire emio_enet2_mdio_mdc,
input  wire emio_enet2_mdio_i,
output wire emio_enet2_mdio_o,
output wire emio_enet2_mdio_t_n,

output wire [2:0] emio_enet3_speed_mode,
input  wire emio_enet3_gmii_crs,
input  wire emio_enet3_gmii_col,
input  wire [7:0] emio_enet3_gmii_rxd,
output wire [7:0] emio_enet3_gmii_txd,
output wire emio_enet3_gmii_tx_en,
output wire emio_enet3_gmii_tx_er,
output wire emio_enet3_mdio_mdc,
input  wire emio_enet3_mdio_i,
output wire emio_enet3_mdio_o,
output wire emio_enet3_mdio_t_n,

input  wire emio_enet0_tx_r_data_rdy,
output wire emio_enet0_tx_r_rd,
input  wire emio_enet0_tx_r_valid,
input  wire [7:0] emio_enet0_tx_r_data,
input  wire emio_enet0_tx_r_sop,
input  wire emio_enet0_tx_r_eop,
input  wire emio_enet0_tx_r_err,
input  wire emio_enet0_tx_r_underflow,
input  wire emio_enet0_tx_r_flushed,
input  wire emio_enet0_tx_r_control,
output wire emio_enet0_dma_tx_end_tog,
input  wire emio_enet0_dma_tx_status_tog,
output wire [3:0] emio_enet0_tx_r_status,
output wire emio_enet0_rx_w_wr,
output wire [7:0] emio_enet0_rx_w_data,
output wire emio_enet0_rx_w_sop,
output wire emio_enet0_rx_w_eop,
output wire [44:0] emio_enet0_rx_w_status,
output wire emio_enet0_rx_w_err,
input  wire emio_enet0_rx_w_overflow,
input  wire emio_enet0_signal_detect,
output wire emio_enet0_rx_w_flush,
output wire emio_enet0_tx_r_fixed_lat,

input  wire emio_enet1_tx_r_data_rdy,
output wire emio_enet1_tx_r_rd,
input  wire emio_enet1_tx_r_valid,
input  wire [7:0] emio_enet1_tx_r_data,
input  wire emio_enet1_tx_r_sop,
input  wire emio_enet1_tx_r_eop,
input  wire emio_enet1_tx_r_err,
input  wire emio_enet1_tx_r_underflow,
input  wire emio_enet1_tx_r_flushed,
input  wire emio_enet1_tx_r_control,
output wire emio_enet1_dma_tx_end_tog,
input  wire emio_enet1_dma_tx_status_tog,
output wire [3:0] emio_enet1_tx_r_status,
output wire emio_enet1_rx_w_wr,
output wire [7:0] emio_enet1_rx_w_data,
output wire emio_enet1_rx_w_sop,
output wire emio_enet1_rx_w_eop,
output wire [44:0] emio_enet1_rx_w_status,
output wire emio_enet1_rx_w_err,
input  wire emio_enet1_rx_w_overflow,
input  wire emio_enet1_signal_detect,
output wire emio_enet1_rx_w_flush,
output wire emio_enet1_tx_r_fixed_lat,

input  wire emio_enet2_tx_r_data_rdy,
output wire emio_enet2_tx_r_rd,
input  wire emio_enet2_tx_r_valid,
input  wire [7:0] emio_enet2_tx_r_data,
input  wire emio_enet2_tx_r_sop,
input  wire emio_enet2_tx_r_eop,
input  wire emio_enet2_tx_r_err,
input  wire emio_enet2_tx_r_underflow,
input  wire emio_enet2_tx_r_flushed,
input  wire emio_enet2_tx_r_control,
output wire emio_enet2_dma_tx_end_tog,
input  wire emio_enet2_dma_tx_status_tog,
output wire [3:0] emio_enet2_tx_r_status,
output wire emio_enet2_rx_w_wr,
output wire [7:0] emio_enet2_rx_w_data,
output wire emio_enet2_rx_w_sop,
output wire emio_enet2_rx_w_eop,
output wire [44:0] emio_enet2_rx_w_status,
output wire emio_enet2_rx_w_err,
input  wire emio_enet2_rx_w_overflow,
input  wire emio_enet2_signal_detect,
output wire emio_enet2_rx_w_flush,
output wire emio_enet2_tx_r_fixed_lat,

input  wire emio_enet3_tx_r_data_rdy,
output wire emio_enet3_tx_r_rd,
input  wire emio_enet3_tx_r_valid,
input  wire [7:0] emio_enet3_tx_r_data,
input  wire emio_enet3_tx_r_sop,
input  wire emio_enet3_tx_r_eop,
input  wire emio_enet3_tx_r_err,
input  wire emio_enet3_tx_r_underflow,
input  wire emio_enet3_tx_r_flushed,
input  wire emio_enet3_tx_r_control,
output wire emio_enet3_dma_tx_end_tog,
input  wire emio_enet3_dma_tx_status_tog,
output wire [3:0] emio_enet3_tx_r_status,
output wire emio_enet3_rx_w_wr,
output wire [7:0] emio_enet3_rx_w_data,
output wire emio_enet3_rx_w_sop,
output wire emio_enet3_rx_w_eop,
output wire [44:0] emio_enet3_rx_w_status,
output wire emio_enet3_rx_w_err,
input  wire emio_enet3_rx_w_overflow,
input  wire emio_enet3_signal_detect,
output wire emio_enet3_rx_w_flush,
output wire emio_enet3_tx_r_fixed_lat,

output wire emio_enet0_tx_sof,
output wire emio_enet0_sync_frame_tx,
output wire emio_enet0_delay_req_tx,
output wire emio_enet0_pdelay_req_tx,
output wire emio_enet0_pdelay_resp_tx,
output wire emio_enet0_rx_sof,
output wire emio_enet0_sync_frame_rx,
output wire emio_enet0_delay_req_rx,
output wire emio_enet0_pdelay_req_rx,
output wire emio_enet0_pdelay_resp_rx,
input  wire [1:0] emio_enet0_tsu_inc_ctrl,
output wire emio_enet0_tsu_timer_cmp_val,
output wire emio_enet1_tx_sof,
output wire emio_enet1_sync_frame_tx,
output wire emio_enet1_delay_req_tx,
output wire emio_enet1_pdelay_req_tx,
output wire emio_enet1_pdelay_resp_tx,
output wire emio_enet1_rx_sof,
output wire emio_enet1_sync_frame_rx,
output wire emio_enet1_delay_req_rx,
output wire emio_enet1_pdelay_req_rx,
output wire emio_enet1_pdelay_resp_rx,
input  wire [1:0] emio_enet1_tsu_inc_ctrl,
output wire emio_enet1_tsu_timer_cmp_val,
output wire emio_enet2_tx_sof,
output wire emio_enet2_sync_frame_tx,
output wire emio_enet2_delay_req_tx,
output wire emio_enet2_pdelay_req_tx,
output wire emio_enet2_pdelay_resp_tx,
output wire emio_enet2_rx_sof,
output wire emio_enet2_sync_frame_rx,
output wire emio_enet2_delay_req_rx,
output wire emio_enet2_pdelay_req_rx,
output wire emio_enet2_pdelay_resp_rx,
input  wire [1:0] emio_enet2_tsu_inc_ctrl,
output wire emio_enet2_tsu_timer_cmp_val,
output wire emio_enet3_tx_sof,
output wire emio_enet3_sync_frame_tx,
output wire emio_enet3_delay_req_tx,
output wire emio_enet3_pdelay_req_tx,
output wire emio_enet3_pdelay_resp_tx,
output wire emio_enet3_rx_sof,
output wire emio_enet3_sync_frame_rx,
output wire emio_enet3_delay_req_rx,
output wire emio_enet3_pdelay_req_rx,
output wire emio_enet3_pdelay_resp_rx,
input  wire [1:0] emio_enet3_tsu_inc_ctrl,
output wire emio_enet3_tsu_timer_cmp_val,

input  wire emio_enet3_gmii_rx_er,
input  wire emio_enet3_gmii_rx_dv,
output wire [93:0] emio_enet0_enet_tsu_timer_cnt,
input  wire emio_enet0_ext_int_in,
input  wire emio_enet1_ext_int_in,
input  wire emio_enet2_ext_int_in,
input  wire emio_enet3_ext_int_in,
output wire [1:0] emio_enet0_dma_bus_width,
output wire [1:0] emio_enet1_dma_bus_width,
output wire [1:0] emio_enet2_dma_bus_width,
output wire [1:0] emio_enet3_dma_bus_width,

input  wire [95:0] emio_gpio_i,
output wire [95:0] emio_gpio_o,
output wire [95:0] emio_gpio_t_n,

input  wire emio_i2c0_scl_i,
output wire emio_i2c0_scl_o,
output wire emio_i2c0_scl_t_n,
input  wire emio_i2c0_sda_i,
output wire emio_i2c0_sda_o,
output wire emio_i2c0_sda_t_n,

input  wire emio_i2c1_scl_i,
output wire emio_i2c1_scl_o,
output wire emio_i2c1_scl_t_n,
input  wire emio_i2c1_sda_i,
output wire emio_i2c1_sda_o,
output wire emio_i2c1_sda_t_n,

output wire emio_uart0_txd,
input  wire emio_uart0_rxd,
input  wire emio_uart0_ctsn,
output wire emio_uart0_rtsn,
input  wire emio_uart0_dsrn,
input  wire emio_uart0_dcdn,
input  wire emio_uart0_rin,
output wire emio_uart0_dtrn,

output wire emio_uart1_txd,
input  wire emio_uart1_rxd,
input  wire emio_uart1_ctsn,
output wire emio_uart1_rtsn,
input  wire emio_uart1_dsrn,
input  wire emio_uart1_dcdn,
input  wire emio_uart1_rin,
output wire emio_uart1_dtrn,

output wire emio_sdio0_cmdout,
input  wire emio_sdio0_cmdin,
output wire emio_sdio0_cmdena_n,
input  wire [7:0] emio_sdio0_datain,
output wire [7:0] emio_sdio0_dataout,
output wire [7:0] emio_sdio0_dataena_n,
input  wire emio_sdio0_cd_n,
input  wire emio_sdio0_wp,
output wire emio_sdio0_ledcontrol,
output wire emio_sdio0_buspower,
output wire [2:0] emio_sdio0_bus_volt,

output wire emio_sdio1_cmdout,
input  wire emio_sdio1_cmdin,
output wire emio_sdio1_cmdena_n,
input  wire [7:0] emio_sdio1_datain,
output wire [7:0] emio_sdio1_dataout,
output wire [7:0] emio_sdio1_dataena_n,
input  wire emio_sdio1_cd_n,
input  wire emio_sdio1_wp,
output wire emio_sdio1_ledcontrol,
output wire emio_sdio1_buspower,
output wire [2:0] emio_sdio1_bus_volt,

input  wire emio_spi0_m_i,
output wire emio_spi0_m_o,
output wire emio_spi0_mo_t_n,
input  wire emio_spi0_s_i,
output wire emio_spi0_s_o,
output wire emio_spi0_so_t_n,
input  wire emio_spi0_ss_i_n,
output wire emio_spi0_ss_o_n,
output wire emio_spi0_ss1_o_n,
output wire emio_spi0_ss2_o_n,
output wire emio_spi0_ss_n_t_n,
input  wire emio_spi0_sclk_i,
output wire emio_spi0_sclk_o,
output wire emio_spi0_sclk_t_n,

input  wire emio_spi1_m_i,
output wire emio_spi1_m_o,
output wire emio_spi1_mo_t_n,
input  wire emio_spi1_s_i,
output wire emio_spi1_s_o,
output wire emio_spi1_so_t_n,
input  wire emio_spi1_ss_i_n,
output wire emio_spi1_ss_o_n,
output wire emio_spi1_ss1_o_n,
output wire emio_spi1_ss2_o_n,
output wire emio_spi1_ss_n_t_n,
input  wire emio_spi1_sclk_i,
output wire emio_spi1_sclk_o,
output wire emio_spi1_sclk_t_n,

output wire ps_pl_tracectl,
output wire [31:0] ps_pl_tracedata,

output wire [2:0] emio_ttc0_wave_o,
output wire [2:0] emio_ttc1_wave_o,
output wire [2:0] emio_ttc2_wave_o,
output wire [2:0] emio_ttc3_wave_o,

output wire emio_wdt0_rst_o,
output wire emio_wdt1_rst_o,

input  wire emio_hub_port_overcrnt_usb3_0,
input  wire emio_hub_port_overcrnt_usb3_1,
input  wire emio_hub_port_overcrnt_usb2_0,
input  wire emio_hub_port_overcrnt_usb2_1,
output wire emio_u2dsport_vbus_ctrl_usb3_0,
output wire emio_u2dsport_vbus_ctrl_usb3_1,
output wire emio_u3dsport_vbus_ctrl_usb3_0,
output wire emio_u3dsport_vbus_ctrl_usb3_1,

input  wire [7:0] pl2adma_cvld,
input  wire [7:0] pl2adma_tack,
output wire [7:0] adma2pl_cack,
output wire [7:0] adma2pl_tvld,

input  wire [7:0] perif_gdma_cvld,
input  wire [7:0] perif_gdma_tack,
output wire [7:0] gdma_perif_cack,
output wire [7:0] gdma_perif_tvld,

input  wire [3:0] pl_clock_stop,

input  wire dp_live_video_in_vsync,
input  wire dp_live_video_in_hsync,
input  wire dp_live_video_in_de,
input  wire [35:0] dp_live_video_in_pixel1,
output wire dp_video_out_hsync,
output wire dp_video_out_vsync,
output wire [35:0] dp_video_out_pixel1,
input  wire dp_aux_data_in,
output wire dp_aux_data_out,
output wire dp_aux_data_oe_n,
input  wire [7:0] dp_live_gfx_alpha_in,
input  wire [35:0] dp_live_gfx_pixel1_in,
input  wire dp_hot_plug_detect,
input  wire dp_external_custom_event1,
input  wire dp_external_custom_event2,
input  wire dp_external_vsync_event,
output wire dp_live_video_de_out,

input  wire pl_ps_eventi,
output wire ps_pl_evento,
output wire [3:0] ps_pl_standbywfe,
output wire [3:0] ps_pl_standbywfi,
input  wire [3:0] pl_ps_apugic_irq,
input  wire [3:0] pl_ps_apugic_fiq,

input  wire rpu_eventi0,
input  wire rpu_eventi1,
output wire rpu_evento0,
output wire rpu_evento1,
input  wire nfiq0_lpd_rpu,
input  wire nfiq1_lpd_rpu,
input  wire nirq0_lpd_rpu,
input  wire nirq1_lpd_rpu,

output wire irq_ipi_pl_0,
output wire irq_ipi_pl_1,
output wire irq_ipi_pl_2,
output wire irq_ipi_pl_3,

input  wire [59:0] stm_event,

// ftm
input  wire [3:0] pl_ps_trigack,
input  wire [3:0] pl_ps_trigger,
output wire [3:0] ps_pl_trigack,
output wire [3:0] ps_pl_trigger,
output wire [31:0] ftm_gpo,
input  wire [31:0] ftm_gpi,

input  wire [7:0] pl_ps_irq0,
input  wire [7:0] pl_ps_irq1,

output wire ps_to_pl_reset0_n,
output wire ps_to_pl_reset1_n,
output wire ps_to_pl_reset2_n,
output wire ps_to_pl_reset3_n,

output wire ps_to_pl_irq_can0,
output wire ps_to_pl_irq_can1,
output wire ps_to_pl_irq_enet0,
output wire ps_to_pl_irq_enet1,
output wire ps_to_pl_irq_enet2,
output wire ps_to_pl_irq_enet3,
output wire ps_to_pl_irq_enet0_wake,
output wire ps_to_pl_irq_enet1_wake,
output wire ps_to_pl_irq_enet2_wake,
output wire ps_to_pl_irq_enet3_wake,
output wire ps_to_pl_irq_gpio,
output wire ps_to_pl_irq_i2c0,
output wire ps_to_pl_irq_i2c1,
output wire ps_to_pl_irq_uart0,
output wire ps_to_pl_irq_uart1,
output wire ps_to_pl_irq_sdio0,
output wire ps_to_pl_irq_sdio1,
output wire ps_to_pl_irq_sdio0_wake,
output wire ps_to_pl_irq_sdio1_wake,
output wire ps_to_pl_irq_spi0,
output wire ps_to_pl_irq_spi1,
output wire ps_to_pl_irq_qspi,
output wire ps_to_pl_irq_ttc0_0,
output wire ps_to_pl_irq_ttc0_1,
output wire ps_to_pl_irq_ttc0_2,
output wire ps_to_pl_irq_ttc1_0,
output wire ps_to_pl_irq_ttc1_1,
output wire ps_to_pl_irq_ttc1_2,
output wire ps_to_pl_irq_ttc2_0,
output wire ps_to_pl_irq_ttc2_1,
output wire ps_to_pl_irq_ttc2_2,
output wire ps_to_pl_irq_ttc3_0,
output wire ps_to_pl_irq_ttc3_1,
output wire ps_to_pl_irq_ttc3_2,
output wire ps_to_pl_irq_csu_pmu_wdt,
output wire ps_to_pl_irq_lp_wdt,
output wire [3:0] ps_to_pl_irq_usb3_0_endpoint,
output wire ps_to_pl_irq_usb3_0_otg,
output wire [3:0] ps_to_pl_irq_usb3_1_endpoint,
output wire ps_to_pl_irq_usb3_1_otg,
output wire [7:0] ps_to_pl_irq_adma_chan,
output wire [1:0] ps_to_pl_irq_usb3_0_pmu_wakeup,
output wire [7:0] ps_to_pl_irq_gdma_chan,
output wire ps_to_pl_irq_csu,
output wire ps_to_pl_irq_csu_dma,
output wire ps_to_pl_irq_efuse,
output wire ps_to_pl_irq_xmpu_lpd,
output wire ps_to_pl_irq_ddr_ss,
output wire ps_to_pl_irq_nand,
output wire ps_to_pl_irq_fp_wdt,
output wire [1:0] ps_to_pl_irq_pcie_msi,
output wire ps_to_pl_irq_pcie_legacy,
output wire ps_to_pl_irq_pcie_dma,
output wire ps_to_pl_irq_pcie_msc,
output wire ps_to_pl_irq_dport,
output wire ps_to_pl_irq_fpd_apb_int,
output wire ps_to_pl_irq_fpd_atb_error,
output wire ps_to_pl_irq_dpdma,
output wire ps_to_pl_irq_apm_fpd,
output wire ps_to_pl_irq_gpu,
output wire ps_to_pl_irq_sata,
output wire ps_to_pl_irq_xmpu_fpd,
output wire [3:0] ps_to_pl_irq_apu_cpumnt,
output wire [3:0] ps_to_pl_irq_apu_cti,
output wire [3:0] ps_to_pl_irq_apu_pmu,
output wire [3:0] ps_to_pl_irq_apu_comm,
output wire ps_to_pl_irq_apu_l2err,
output wire ps_to_pl_irq_apu_exterr,
output wire ps_to_pl_irq_apu_regs,
output wire ps_to_pl_irq_intf_ppd_cci,
output wire ps_to_pl_irq_intf_fpd_smmu,
output wire ps_to_pl_irq_atb_err_lpd,
output wire ps_to_pl_irq_aib_axi,
output wire ps_to_pl_irq_ams,
output wire ps_to_pl_irq_lpd_apm,
output wire ps_to_pl_irq_rtc_alaram,
output wire ps_to_pl_irq_rtc_seconds,
output wire ps_to_pl_irq_clkmon,
output wire ps_to_pl_irq_ipi_channel0,
output wire ps_to_pl_irq_ipi_channel1,
output wire ps_to_pl_irq_ipi_channel2,
output wire ps_to_pl_irq_ipi_channel7,
output wire ps_to_pl_irq_ipi_channel8,
output wire ps_to_pl_irq_ipi_channel9,
output wire ps_to_pl_irq_ipi_channel10,
output wire [1:0] ps_to_pl_irq_rpu_pm,
output wire ps_to_pl_irq_ocm_error,
output wire ps_to_pl_irq_lpd_apb_intr,
output wire ps_to_pl_irq_r5_core0_ecc_error,
output wire ps_to_pl_irq_r5_core1_ecc_error,


output wire osc_rtc_clk,

input  wire [31:0] pl_pmu_gpi,
output wire [31:0] pmu_pl_gpo,
input  wire aib_pmu_afifm_fpd_ack,
input  wire aib_pmu_afifm_lpd_ack,
output wire pmu_aib_afifm_fpd_req,
output wire pmu_aib_afifm_lpd_req,
output wire [46:0] pmu_error_to_pl,
input  wire [3:0] pmu_error_from_pl,

input  wire ddrc_ext_refresh_rank0_req,
input  wire ddrc_ext_refresh_rank1_req,
input  wire pl_acpinact,

input  [31:0] pstp_pl_in,
output [31:0] pstp_pl_out,
input  [31:0] pstp_pl_ts
);

// these are not used sinks for irq lines form PS
wire [18:0] irq_lpd_dev_null;
wire [19:0] irq_fpd_dev_null;

// unclear what these are
wire pss_alto_core_pad_mgttxn0out;
wire pss_alto_core_pad_mgttxp0out;
wire pss_alto_core_pad_mgttxn1out;
wire pss_alto_core_pad_mgttxp1out;
wire pss_alto_core_pad_mgttxn2out;
wire pss_alto_core_pad_mgttxp2out;
wire pss_alto_core_pad_mgttxn3out;
wire pss_alto_core_pad_mgttxp3out;
wire pss_alto_core_pad_pado;

// rename the gpio reset lins
assign ps_to_pl_reset0_n = emio_gpio_i[95];
assign ps_to_pl_reset1_n = emio_gpio_i[94];
assign ps_to_pl_reset2_n = emio_gpio_i[93];
assign ps_to_pl_reset3_n = emio_gpio_i[92];

PS8 PS8_i  (
.MAXIGP0ACLK (clk_ps_to_pl_axi_hpm0_fpd),
.MAXIGP0AWID (ps_to_pl_axi_hpm0_fpd_awid),
.MAXIGP0AWADDR (ps_to_pl_axi_hpm0_fpd_awaddr),
.MAXIGP0AWLEN (ps_to_pl_axi_hpm0_fpd_awlen),
.MAXIGP0AWSIZE (ps_to_pl_axi_hpm0_fpd_awsize),
.MAXIGP0AWBURST (ps_to_pl_axi_hpm0_fpd_awburst),
.MAXIGP0AWLOCK (ps_to_pl_axi_hpm0_fpd_awlock),
.MAXIGP0AWCACHE (ps_to_pl_axi_hpm0_fpd_awcache),
.MAXIGP0AWPROT (ps_to_pl_axi_hpm0_fpd_awprot),
.MAXIGP0AWVALID (ps_to_pl_axi_hpm0_fpd_awvalid),
.MAXIGP0AWUSER (ps_to_pl_axi_hpm0_fpd_awuser),
.MAXIGP0AWREADY (ps_to_pl_axi_hpm0_fpd_awready),
.MAXIGP0WDATA (ps_to_pl_axi_hpm0_fpd_wdata),
.MAXIGP0WSTRB (ps_to_pl_axi_hpm0_fpd_wstrb),
.MAXIGP0WLAST (ps_to_pl_axi_hpm0_fpd_wlast),
.MAXIGP0WVALID (ps_to_pl_axi_hpm0_fpd_wvalid),
.MAXIGP0WREADY (ps_to_pl_axi_hpm0_fpd_wready),
.MAXIGP0BID (ps_to_pl_axi_hpm0_fpd_bid),
.MAXIGP0BRESP (ps_to_pl_axi_hpm0_fpd_bresp),
.MAXIGP0BVALID (ps_to_pl_axi_hpm0_fpd_bvalid),
.MAXIGP0BREADY (ps_to_pl_axi_hpm0_fpd_bready),
.MAXIGP0ARID (ps_to_pl_axi_hpm0_fpd_arid),
.MAXIGP0ARADDR (ps_to_pl_axi_hpm0_fpd_araddr),
.MAXIGP0ARLEN (ps_to_pl_axi_hpm0_fpd_arlen),
.MAXIGP0ARSIZE (ps_to_pl_axi_hpm0_fpd_arsize),
.MAXIGP0ARBURST (ps_to_pl_axi_hpm0_fpd_arburst),
.MAXIGP0ARLOCK (ps_to_pl_axi_hpm0_fpd_arlock),
.MAXIGP0ARCACHE (ps_to_pl_axi_hpm0_fpd_arcache),
.MAXIGP0ARPROT (ps_to_pl_axi_hpm0_fpd_arprot),
.MAXIGP0ARVALID (ps_to_pl_axi_hpm0_fpd_arvalid),
.MAXIGP0ARUSER (ps_to_pl_axi_hpm0_fpd_aruser),
.MAXIGP0ARREADY (ps_to_pl_axi_hpm0_fpd_arready),
.MAXIGP0RID (ps_to_pl_axi_hpm0_fpd_rid),
.MAXIGP0RDATA (ps_to_pl_axi_hpm0_fpd_rdata),
.MAXIGP0RRESP (ps_to_pl_axi_hpm0_fpd_rresp),
.MAXIGP0RLAST (ps_to_pl_axi_hpm0_fpd_rlast),
.MAXIGP0RVALID (ps_to_pl_axi_hpm0_fpd_rvalid),
.MAXIGP0RREADY (ps_to_pl_axi_hpm0_fpd_rready),
.MAXIGP0AWQOS (ps_to_pl_axi_hpm0_fpd_awqos),
.MAXIGP0ARQOS (ps_to_pl_axi_hpm0_fpd_arqos),
.MAXIGP1ACLK (clk_ps_to_pl_axi_hpm1_fpd),
.MAXIGP1AWID (ps_to_pl_axi_hpm1_fpd_awid),
.MAXIGP1AWADDR (ps_to_pl_axi_hpm1_fpd_awaddr),
.MAXIGP1AWLEN (ps_to_pl_axi_hpm1_fpd_awlen),
.MAXIGP1AWSIZE (ps_to_pl_axi_hpm1_fpd_awsize),
.MAXIGP1AWBURST (ps_to_pl_axi_hpm1_fpd_awburst),
.MAXIGP1AWLOCK (ps_to_pl_axi_hpm1_fpd_awlock),
.MAXIGP1AWCACHE (ps_to_pl_axi_hpm1_fpd_awcache),
.MAXIGP1AWPROT (ps_to_pl_axi_hpm1_fpd_awprot),
.MAXIGP1AWVALID (ps_to_pl_axi_hpm1_fpd_awvalid),
.MAXIGP1AWUSER (ps_to_pl_axi_hpm1_fpd_awuser),
.MAXIGP1AWREADY (ps_to_pl_axi_hpm1_fpd_awready),
.MAXIGP1WDATA (ps_to_pl_axi_hpm1_fpd_wdata),
.MAXIGP1WSTRB (ps_to_pl_axi_hpm1_fpd_wstrb),
.MAXIGP1WLAST (ps_to_pl_axi_hpm1_fpd_wlast),
.MAXIGP1WVALID (ps_to_pl_axi_hpm1_fpd_wvalid),
.MAXIGP1WREADY (ps_to_pl_axi_hpm1_fpd_wready),
.MAXIGP1BID (ps_to_pl_axi_hpm1_fpd_bid),
.MAXIGP1BRESP (ps_to_pl_axi_hpm1_fpd_bresp),
.MAXIGP1BVALID (ps_to_pl_axi_hpm1_fpd_bvalid),
.MAXIGP1BREADY (ps_to_pl_axi_hpm1_fpd_bready),
.MAXIGP1ARID (ps_to_pl_axi_hpm1_fpd_arid),
.MAXIGP1ARADDR (ps_to_pl_axi_hpm1_fpd_araddr),
.MAXIGP1ARLEN (ps_to_pl_axi_hpm1_fpd_arlen),
.MAXIGP1ARSIZE (ps_to_pl_axi_hpm1_fpd_arsize),
.MAXIGP1ARBURST (ps_to_pl_axi_hpm1_fpd_arburst),
.MAXIGP1ARLOCK (ps_to_pl_axi_hpm1_fpd_arlock),
.MAXIGP1ARCACHE (ps_to_pl_axi_hpm1_fpd_arcache),
.MAXIGP1ARPROT (ps_to_pl_axi_hpm1_fpd_arprot),
.MAXIGP1ARVALID (ps_to_pl_axi_hpm1_fpd_arvalid),
.MAXIGP1ARUSER (ps_to_pl_axi_hpm1_fpd_aruser),
.MAXIGP1ARREADY (ps_to_pl_axi_hpm1_fpd_arready),
.MAXIGP1RID (ps_to_pl_axi_hpm1_fpd_rid),
.MAXIGP1RDATA (ps_to_pl_axi_hpm1_fpd_rdata),
.MAXIGP1RRESP (ps_to_pl_axi_hpm1_fpd_rresp),
.MAXIGP1RLAST (ps_to_pl_axi_hpm1_fpd_rlast),
.MAXIGP1RVALID (ps_to_pl_axi_hpm1_fpd_rvalid),
.MAXIGP1RREADY (ps_to_pl_axi_hpm1_fpd_rready),
.MAXIGP1AWQOS (ps_to_pl_axi_hpm1_fpd_awqos),
.MAXIGP1ARQOS (ps_to_pl_axi_hpm1_fpd_arqos),
.MAXIGP2ACLK (clk_ps_to_pl_axi_hpm0_lpd),
.MAXIGP2AWID (ps_to_pl_axi_hpm0_lpd_awid),
.MAXIGP2AWADDR (ps_to_pl_axi_hpm0_lpd_awaddr),
.MAXIGP2AWLEN (ps_to_pl_axi_hpm0_lpd_awlen),
.MAXIGP2AWSIZE (ps_to_pl_axi_hpm0_lpd_awsize),
.MAXIGP2AWBURST (ps_to_pl_axi_hpm0_lpd_awburst),
.MAXIGP2AWLOCK (ps_to_pl_axi_hpm0_lpd_awlock),
.MAXIGP2AWCACHE (ps_to_pl_axi_hpm0_lpd_awcache),
.MAXIGP2AWPROT (ps_to_pl_axi_hpm0_lpd_awprot),
.MAXIGP2AWVALID (ps_to_pl_axi_hpm0_lpd_awvalid),
.MAXIGP2AWUSER (ps_to_pl_axi_hpm0_lpd_awuser),
.MAXIGP2AWREADY (ps_to_pl_axi_hpm0_lpd_awready),
.MAXIGP2WDATA (ps_to_pl_axi_hpm0_lpd_wdata),
.MAXIGP2WSTRB (ps_to_pl_axi_hpm0_lpd_wstrb),
.MAXIGP2WLAST (ps_to_pl_axi_hpm0_lpd_wlast),
.MAXIGP2WVALID (ps_to_pl_axi_hpm0_lpd_wvalid),
.MAXIGP2WREADY (ps_to_pl_axi_hpm0_lpd_wready),
.MAXIGP2BID (ps_to_pl_axi_hpm0_lpd_bid),
.MAXIGP2BRESP (ps_to_pl_axi_hpm0_lpd_bresp),
.MAXIGP2BVALID (ps_to_pl_axi_hpm0_lpd_bvalid),
.MAXIGP2BREADY (ps_to_pl_axi_hpm0_lpd_bready),
.MAXIGP2ARID (ps_to_pl_axi_hpm0_lpd_arid),
.MAXIGP2ARADDR (ps_to_pl_axi_hpm0_lpd_araddr),
.MAXIGP2ARLEN (ps_to_pl_axi_hpm0_lpd_arlen),
.MAXIGP2ARSIZE (ps_to_pl_axi_hpm0_lpd_arsize),
.MAXIGP2ARBURST (ps_to_pl_axi_hpm0_lpd_arburst),
.MAXIGP2ARLOCK (ps_to_pl_axi_hpm0_lpd_arlock),
.MAXIGP2ARCACHE (ps_to_pl_axi_hpm0_lpd_arcache),
.MAXIGP2ARPROT (ps_to_pl_axi_hpm0_lpd_arprot),
.MAXIGP2ARVALID (ps_to_pl_axi_hpm0_lpd_arvalid),
.MAXIGP2ARUSER (ps_to_pl_axi_hpm0_lpd_aruser),
.MAXIGP2ARREADY (ps_to_pl_axi_hpm0_lpd_arready),
.MAXIGP2RID (ps_to_pl_axi_hpm0_lpd_rid),
.MAXIGP2RDATA (ps_to_pl_axi_hpm0_lpd_rdata),
.MAXIGP2RRESP (ps_to_pl_axi_hpm0_lpd_rresp),
.MAXIGP2RLAST (ps_to_pl_axi_hpm0_lpd_rlast),
.MAXIGP2RVALID (ps_to_pl_axi_hpm0_lpd_rvalid),
.MAXIGP2RREADY (ps_to_pl_axi_hpm0_lpd_rready),
.MAXIGP2AWQOS (ps_to_pl_axi_hpm0_lpd_awqos),
.MAXIGP2ARQOS (ps_to_pl_axi_hpm0_lpd_arqos),
.SAXIGP0RCLK (clk_pl_to_ps_axi_hpc0_fpd_read),
.SAXIGP0WCLK (clk_pl_to_ps_axi_hpc0_fpd_write),
.SAXIGP0ARUSER (pl_to_ps_axi_hpc0_fpd_aruser),
.SAXIGP0AWUSER (pl_to_ps_axi_hpc0_fpd_awuser),
.SAXIGP0AWID (pl_to_ps_axi_hpc0_fpd_awid),
.SAXIGP0AWADDR (pl_to_ps_axi_hpc0_fpd_awaddr),
.SAXIGP0AWLEN (pl_to_ps_axi_hpc0_fpd_awlen),
.SAXIGP0AWSIZE (pl_to_ps_axi_hpc0_fpd_awsize),
.SAXIGP0AWBURST (pl_to_ps_axi_hpc0_fpd_awburst),
.SAXIGP0AWLOCK (pl_to_ps_axi_hpc0_fpd_awlock),
.SAXIGP0AWCACHE (pl_to_ps_axi_hpc0_fpd_awcache),
.SAXIGP0AWPROT (pl_to_ps_axi_hpc0_fpd_awprot),
.SAXIGP0AWVALID (pl_to_ps_axi_hpc0_fpd_awvalid),
.SAXIGP0AWREADY (pl_to_ps_axi_hpc0_fpd_awready),
.SAXIGP0WDATA (pl_to_ps_axi_hpc0_fpd_wdata),
.SAXIGP0WSTRB (pl_to_ps_axi_hpc0_fpd_wstrb),
.SAXIGP0WLAST (pl_to_ps_axi_hpc0_fpd_wlast),
.SAXIGP0WVALID (pl_to_ps_axi_hpc0_fpd_wvalid),
.SAXIGP0WREADY (pl_to_ps_axi_hpc0_fpd_wready),
.SAXIGP0BID (pl_to_ps_axi_hpc0_fpd_bid),
.SAXIGP0BRESP (pl_to_ps_axi_hpc0_fpd_bresp),
.SAXIGP0BVALID (pl_to_ps_axi_hpc0_fpd_bvalid),
.SAXIGP0BREADY (pl_to_ps_axi_hpc0_fpd_bready),
.SAXIGP0ARID (pl_to_ps_axi_hpc0_fpd_arid),
.SAXIGP0ARADDR (pl_to_ps_axi_hpc0_fpd_araddr),
.SAXIGP0ARLEN (pl_to_ps_axi_hpc0_fpd_arlen),
.SAXIGP0ARSIZE (pl_to_ps_axi_hpc0_fpd_arsize),
.SAXIGP0ARBURST (pl_to_ps_axi_hpc0_fpd_arburst),
.SAXIGP0ARLOCK (pl_to_ps_axi_hpc0_fpd_arlock),
.SAXIGP0ARCACHE (pl_to_ps_axi_hpc0_fpd_arcache),
.SAXIGP0ARPROT (pl_to_ps_axi_hpc0_fpd_arprot),
.SAXIGP0ARVALID (pl_to_ps_axi_hpc0_fpd_arvalid),
.SAXIGP0ARREADY (pl_to_ps_axi_hpc0_fpd_arready),
.SAXIGP0RID (pl_to_ps_axi_hpc0_fpd_rid),
.SAXIGP0RDATA (pl_to_ps_axi_hpc0_fpd_rdata),
.SAXIGP0RRESP (pl_to_ps_axi_hpc0_fpd_rresp),
.SAXIGP0RLAST (pl_to_ps_axi_hpc0_fpd_rlast),
.SAXIGP0RVALID (pl_to_ps_axi_hpc0_fpd_rvalid),
.SAXIGP0RREADY (pl_to_ps_axi_hpc0_fpd_rready),
.SAXIGP0AWQOS (pl_to_ps_axi_hpc0_fpd_awqos),
.SAXIGP0ARQOS (pl_to_ps_axi_hpc0_fpd_arqos),
.SAXIGP0RCOUNT (pl_to_ps_axi_hpc0_fpd_rcount),
.SAXIGP0WCOUNT (pl_to_ps_axi_hpc0_fpd_wcount),
.SAXIGP0RACOUNT (pl_to_ps_axi_hpc0_fpd_racount),
.SAXIGP0WACOUNT (pl_to_ps_axi_hpc0_fpd_wacount),
.SAXIGP1RCLK (clk_pl_to_ps_axi_hpc1_fpd_read),
.SAXIGP1WCLK (clk_pl_to_ps_axi_hpc1_fpd_write),
.SAXIGP1ARUSER (pl_to_ps_axi_hpc1_fpd_aruser),
.SAXIGP1AWUSER (pl_to_ps_axi_hpc1_fpd_awuser),
.SAXIGP1AWID (pl_to_ps_axi_hpc1_fpd_awid),
.SAXIGP1AWADDR (pl_to_ps_axi_hpc1_fpd_awaddr),
.SAXIGP1AWLEN (pl_to_ps_axi_hpc1_fpd_awlen),
.SAXIGP1AWSIZE (pl_to_ps_axi_hpc1_fpd_awsize),
.SAXIGP1AWBURST (pl_to_ps_axi_hpc1_fpd_awburst),
.SAXIGP1AWLOCK (pl_to_ps_axi_hpc1_fpd_awlock),
.SAXIGP1AWCACHE (pl_to_ps_axi_hpc1_fpd_awcache),
.SAXIGP1AWPROT (pl_to_ps_axi_hpc1_fpd_awprot),
.SAXIGP1AWVALID (pl_to_ps_axi_hpc1_fpd_awvalid),
.SAXIGP1AWREADY (pl_to_ps_axi_hpc1_fpd_awready),
.SAXIGP1WDATA (pl_to_ps_axi_hpc1_fpd_wdata),
.SAXIGP1WSTRB (pl_to_ps_axi_hpc1_fpd_wstrb),
.SAXIGP1WLAST (pl_to_ps_axi_hpc1_fpd_wlast),
.SAXIGP1WVALID (pl_to_ps_axi_hpc1_fpd_wvalid),
.SAXIGP1WREADY (pl_to_ps_axi_hpc1_fpd_wready),
.SAXIGP1BID (pl_to_ps_axi_hpc1_fpd_bid),
.SAXIGP1BRESP (pl_to_ps_axi_hpc1_fpd_bresp),
.SAXIGP1BVALID (pl_to_ps_axi_hpc1_fpd_bvalid),
.SAXIGP1BREADY (pl_to_ps_axi_hpc1_fpd_bready),
.SAXIGP1ARID (pl_to_ps_axi_hpc1_fpd_arid),
.SAXIGP1ARADDR (pl_to_ps_axi_hpc1_fpd_araddr),
.SAXIGP1ARLEN (pl_to_ps_axi_hpc1_fpd_arlen),
.SAXIGP1ARSIZE (pl_to_ps_axi_hpc1_fpd_arsize),
.SAXIGP1ARBURST (pl_to_ps_axi_hpc1_fpd_arburst),
.SAXIGP1ARLOCK (pl_to_ps_axi_hpc1_fpd_arlock),
.SAXIGP1ARCACHE (pl_to_ps_axi_hpc1_fpd_arcache),
.SAXIGP1ARPROT (pl_to_ps_axi_hpc1_fpd_arprot),
.SAXIGP1ARVALID (pl_to_ps_axi_hpc1_fpd_arvalid),
.SAXIGP1ARREADY (pl_to_ps_axi_hpc1_fpd_arready),
.SAXIGP1RID (pl_to_ps_axi_hpc1_fpd_rid),
.SAXIGP1RDATA (pl_to_ps_axi_hpc1_fpd_rdata),
.SAXIGP1RRESP (pl_to_ps_axi_hpc1_fpd_rresp),
.SAXIGP1RLAST (pl_to_ps_axi_hpc1_fpd_rlast),
.SAXIGP1RVALID (pl_to_ps_axi_hpc1_fpd_rvalid),
.SAXIGP1RREADY (pl_to_ps_axi_hpc1_fpd_rready),
.SAXIGP1AWQOS (pl_to_ps_axi_hpc1_fpd_awqos),
.SAXIGP1ARQOS (pl_to_ps_axi_hpc1_fpd_arqos),
.SAXIGP1RCOUNT (pl_to_ps_axi_hpc1_fpd_rcount),
.SAXIGP1WCOUNT (pl_to_ps_axi_hpc1_fpd_wcount),
.SAXIGP1RACOUNT (pl_to_ps_axi_hpc1_fpd_racount),
.SAXIGP1WACOUNT (pl_to_ps_axi_hpc1_fpd_wacount),
.SAXIGP2RCLK (clk_pl_to_ps_axi_hp0_fpd_read),
.SAXIGP2WCLK (clk_pl_to_ps_axi_hp0_fpd_write),
.SAXIGP2ARUSER (pl_to_ps_axi_hp0_fpd_aruser),
.SAXIGP2AWUSER (pl_to_ps_axi_hp0_fpd_awuser),
.SAXIGP2AWID (pl_to_ps_axi_hp0_fpd_awid),
.SAXIGP2AWADDR (pl_to_ps_axi_hp0_fpd_awaddr),
.SAXIGP2AWLEN (pl_to_ps_axi_hp0_fpd_awlen),
.SAXIGP2AWSIZE (pl_to_ps_axi_hp0_fpd_awsize),
.SAXIGP2AWBURST (pl_to_ps_axi_hp0_fpd_awburst),
.SAXIGP2AWLOCK (pl_to_ps_axi_hp0_fpd_awlock),
.SAXIGP2AWCACHE (pl_to_ps_axi_hp0_fpd_awcache),
.SAXIGP2AWPROT (pl_to_ps_axi_hp0_fpd_awprot),
.SAXIGP2AWVALID (pl_to_ps_axi_hp0_fpd_awvalid),
.SAXIGP2AWREADY (pl_to_ps_axi_hp0_fpd_awready),
.SAXIGP2WDATA (pl_to_ps_axi_hp0_fpd_wdata),
.SAXIGP2WSTRB (pl_to_ps_axi_hp0_fpd_wstrb),
.SAXIGP2WLAST (pl_to_ps_axi_hp0_fpd_wlast),
.SAXIGP2WVALID (pl_to_ps_axi_hp0_fpd_wvalid),
.SAXIGP2WREADY (pl_to_ps_axi_hp0_fpd_wready),
.SAXIGP2BID (pl_to_ps_axi_hp0_fpd_bid),
.SAXIGP2BRESP (pl_to_ps_axi_hp0_fpd_bresp),
.SAXIGP2BVALID (pl_to_ps_axi_hp0_fpd_bvalid),
.SAXIGP2BREADY (pl_to_ps_axi_hp0_fpd_bready),
.SAXIGP2ARID (pl_to_ps_axi_hp0_fpd_arid),
.SAXIGP2ARADDR (pl_to_ps_axi_hp0_fpd_araddr),
.SAXIGP2ARLEN (pl_to_ps_axi_hp0_fpd_arlen),
.SAXIGP2ARSIZE (pl_to_ps_axi_hp0_fpd_arsize),
.SAXIGP2ARBURST (pl_to_ps_axi_hp0_fpd_arburst),
.SAXIGP2ARLOCK (pl_to_ps_axi_hp0_fpd_arlock),
.SAXIGP2ARCACHE (pl_to_ps_axi_hp0_fpd_arcache),
.SAXIGP2ARPROT (pl_to_ps_axi_hp0_fpd_arprot),
.SAXIGP2ARVALID (pl_to_ps_axi_hp0_fpd_arvalid),
.SAXIGP2ARREADY (pl_to_ps_axi_hp0_fpd_arready),
.SAXIGP2RID (pl_to_ps_axi_hp0_fpd_rid),
.SAXIGP2RDATA (pl_to_ps_axi_hp0_fpd_rdata),
.SAXIGP2RRESP (pl_to_ps_axi_hp0_fpd_rresp),
.SAXIGP2RLAST (pl_to_ps_axi_hp0_fpd_rlast),
.SAXIGP2RVALID (pl_to_ps_axi_hp0_fpd_rvalid),
.SAXIGP2RREADY (pl_to_ps_axi_hp0_fpd_rready),
.SAXIGP2AWQOS (pl_to_ps_axi_hp0_fpd_awqos),
.SAXIGP2ARQOS (pl_to_ps_axi_hp0_fpd_arqos),
.SAXIGP2RCOUNT (pl_to_ps_axi_hp0_fpd_rcount),
.SAXIGP2WCOUNT (pl_to_ps_axi_hp0_fpd_wcount),
.SAXIGP2RACOUNT (pl_to_ps_axi_hp0_fpd_racount),
.SAXIGP2WACOUNT (pl_to_ps_axi_hp0_fpd_wacount),
.SAXIGP3RCLK (clk_pl_to_ps_axi_hp1_fpd_read),
.SAXIGP3WCLK (clk_pl_to_ps_axi_hp1_fpd_write),
.SAXIGP3ARUSER (pl_to_ps_axi_hp1_fpd_aruser),
.SAXIGP3AWUSER (pl_to_ps_axi_hp1_fpd_awuser),
.SAXIGP3AWID (pl_to_ps_axi_hp1_fpd_awid),
.SAXIGP3AWADDR (pl_to_ps_axi_hp1_fpd_awaddr),
.SAXIGP3AWLEN (pl_to_ps_axi_hp1_fpd_awlen),
.SAXIGP3AWSIZE (pl_to_ps_axi_hp1_fpd_awsize),
.SAXIGP3AWBURST (pl_to_ps_axi_hp1_fpd_awburst),
.SAXIGP3AWLOCK (pl_to_ps_axi_hp1_fpd_awlock),
.SAXIGP3AWCACHE (pl_to_ps_axi_hp1_fpd_awcache),
.SAXIGP3AWPROT (pl_to_ps_axi_hp1_fpd_awprot),
.SAXIGP3AWVALID (pl_to_ps_axi_hp1_fpd_awvalid),
.SAXIGP3AWREADY (pl_to_ps_axi_hp1_fpd_awready),
.SAXIGP3WDATA (pl_to_ps_axi_hp1_fpd_wdata),
.SAXIGP3WSTRB (pl_to_ps_axi_hp1_fpd_wstrb),
.SAXIGP3WLAST (pl_to_ps_axi_hp1_fpd_wlast),
.SAXIGP3WVALID (pl_to_ps_axi_hp1_fpd_wvalid),
.SAXIGP3WREADY (pl_to_ps_axi_hp1_fpd_wready),
.SAXIGP3BID (pl_to_ps_axi_hp1_fpd_bid),
.SAXIGP3BRESP (pl_to_ps_axi_hp1_fpd_bresp),
.SAXIGP3BVALID (pl_to_ps_axi_hp1_fpd_bvalid),
.SAXIGP3BREADY (pl_to_ps_axi_hp1_fpd_bready),
.SAXIGP3ARID (pl_to_ps_axi_hp1_fpd_arid),
.SAXIGP3ARADDR (pl_to_ps_axi_hp1_fpd_araddr),
.SAXIGP3ARLEN (pl_to_ps_axi_hp1_fpd_arlen),
.SAXIGP3ARSIZE (pl_to_ps_axi_hp1_fpd_arsize),
.SAXIGP3ARBURST (pl_to_ps_axi_hp1_fpd_arburst),
.SAXIGP3ARLOCK (pl_to_ps_axi_hp1_fpd_arlock),
.SAXIGP3ARCACHE (pl_to_ps_axi_hp1_fpd_arcache),
.SAXIGP3ARPROT (pl_to_ps_axi_hp1_fpd_arprot),
.SAXIGP3ARVALID (pl_to_ps_axi_hp1_fpd_arvalid),
.SAXIGP3ARREADY (pl_to_ps_axi_hp1_fpd_arready),
.SAXIGP3RID (pl_to_ps_axi_hp1_fpd_rid),
.SAXIGP3RDATA (pl_to_ps_axi_hp1_fpd_rdata),
.SAXIGP3RRESP (pl_to_ps_axi_hp1_fpd_rresp),
.SAXIGP3RLAST (pl_to_ps_axi_hp1_fpd_rlast),
.SAXIGP3RVALID (pl_to_ps_axi_hp1_fpd_rvalid),
.SAXIGP3RREADY (pl_to_ps_axi_hp1_fpd_rready),
.SAXIGP3AWQOS (pl_to_ps_axi_hp1_fpd_awqos),
.SAXIGP3ARQOS (pl_to_ps_axi_hp1_fpd_arqos),
.SAXIGP3RCOUNT (pl_to_ps_axi_hp1_fpd_rcount),
.SAXIGP3WCOUNT (pl_to_ps_axi_hp1_fpd_wcount),
.SAXIGP3RACOUNT (pl_to_ps_axi_hp1_fpd_racount),
.SAXIGP3WACOUNT (pl_to_ps_axi_hp1_fpd_wacount),
.SAXIGP4RCLK (clk_pl_to_ps_axi_hp2_fpd_read),
.SAXIGP4WCLK (clk_pl_to_ps_axi_hp2_fpd_write),
.SAXIGP4ARUSER (pl_to_ps_axi_hp2_fpd_aruser),
.SAXIGP4AWUSER (pl_to_ps_axi_hp2_fpd_awuser),
.SAXIGP4AWID (pl_to_ps_axi_hp2_fpd_awid),
.SAXIGP4AWADDR (pl_to_ps_axi_hp2_fpd_awaddr),
.SAXIGP4AWLEN (pl_to_ps_axi_hp2_fpd_awlen),
.SAXIGP4AWSIZE (pl_to_ps_axi_hp2_fpd_awsize),
.SAXIGP4AWBURST (pl_to_ps_axi_hp2_fpd_awburst),
.SAXIGP4AWLOCK (pl_to_ps_axi_hp2_fpd_awlock),
.SAXIGP4AWCACHE (pl_to_ps_axi_hp2_fpd_awcache),
.SAXIGP4AWPROT (pl_to_ps_axi_hp2_fpd_awprot),
.SAXIGP4AWVALID (pl_to_ps_axi_hp2_fpd_awvalid),
.SAXIGP4AWREADY (pl_to_ps_axi_hp2_fpd_awready),
.SAXIGP4WDATA (pl_to_ps_axi_hp2_fpd_wdata),
.SAXIGP4WSTRB (pl_to_ps_axi_hp2_fpd_wstrb),
.SAXIGP4WLAST (pl_to_ps_axi_hp2_fpd_wlast),
.SAXIGP4WVALID (pl_to_ps_axi_hp2_fpd_wvalid),
.SAXIGP4WREADY (pl_to_ps_axi_hp2_fpd_wready),
.SAXIGP4BID (pl_to_ps_axi_hp2_fpd_bid),
.SAXIGP4BRESP (pl_to_ps_axi_hp2_fpd_bresp),
.SAXIGP4BVALID (pl_to_ps_axi_hp2_fpd_bvalid),
.SAXIGP4BREADY (pl_to_ps_axi_hp2_fpd_bready),
.SAXIGP4ARID (pl_to_ps_axi_hp2_fpd_arid),
.SAXIGP4ARADDR (pl_to_ps_axi_hp2_fpd_araddr),
.SAXIGP4ARLEN (pl_to_ps_axi_hp2_fpd_arlen),
.SAXIGP4ARSIZE (pl_to_ps_axi_hp2_fpd_arsize),
.SAXIGP4ARBURST (pl_to_ps_axi_hp2_fpd_arburst),
.SAXIGP4ARLOCK (pl_to_ps_axi_hp2_fpd_arlock),
.SAXIGP4ARCACHE (pl_to_ps_axi_hp2_fpd_arcache),
.SAXIGP4ARPROT (pl_to_ps_axi_hp2_fpd_arprot),
.SAXIGP4ARVALID (pl_to_ps_axi_hp2_fpd_arvalid),
.SAXIGP4ARREADY (pl_to_ps_axi_hp2_fpd_arready),
.SAXIGP4RID (pl_to_ps_axi_hp2_fpd_rid),
.SAXIGP4RDATA (pl_to_ps_axi_hp2_fpd_rdata),
.SAXIGP4RRESP (pl_to_ps_axi_hp2_fpd_rresp),
.SAXIGP4RLAST (pl_to_ps_axi_hp2_fpd_rlast),
.SAXIGP4RVALID (pl_to_ps_axi_hp2_fpd_rvalid),
.SAXIGP4RREADY (pl_to_ps_axi_hp2_fpd_rready),
.SAXIGP4AWQOS (pl_to_ps_axi_hp2_fpd_awqos),
.SAXIGP4ARQOS (pl_to_ps_axi_hp2_fpd_arqos),
.SAXIGP4RCOUNT (pl_to_ps_axi_hp2_fpd_rcount),
.SAXIGP4WCOUNT (pl_to_ps_axi_hp2_fpd_wcount),
.SAXIGP4RACOUNT (pl_to_ps_axi_hp2_fpd_racount),
.SAXIGP4WACOUNT (pl_to_ps_axi_hp2_fpd_wacount),
.SAXIGP5RCLK (clk_pl_to_ps_axi_hp3_fpd_read),
.SAXIGP5WCLK (clk_pl_to_ps_axi_hp3_fpd_write),
.SAXIGP5ARUSER (pl_to_ps_axi_hp3_fpd_aruser),
.SAXIGP5AWUSER (pl_to_ps_axi_hp3_fpd_awuser),
.SAXIGP5AWID (pl_to_ps_axi_hp3_fpd_awid),
.SAXIGP5AWADDR (pl_to_ps_axi_hp3_fpd_awaddr),
.SAXIGP5AWLEN (pl_to_ps_axi_hp3_fpd_awlen),
.SAXIGP5AWSIZE (pl_to_ps_axi_hp3_fpd_awsize),
.SAXIGP5AWBURST (pl_to_ps_axi_hp3_fpd_awburst),
.SAXIGP5AWLOCK (pl_to_ps_axi_hp3_fpd_awlock),
.SAXIGP5AWCACHE (pl_to_ps_axi_hp3_fpd_awcache),
.SAXIGP5AWPROT (pl_to_ps_axi_hp3_fpd_awprot),
.SAXIGP5AWVALID (pl_to_ps_axi_hp3_fpd_awvalid),
.SAXIGP5AWREADY (pl_to_ps_axi_hp3_fpd_awready),
.SAXIGP5WDATA (pl_to_ps_axi_hp3_fpd_wdata),
.SAXIGP5WSTRB (pl_to_ps_axi_hp3_fpd_wstrb),
.SAXIGP5WLAST (pl_to_ps_axi_hp3_fpd_wlast),
.SAXIGP5WVALID (pl_to_ps_axi_hp3_fpd_wvalid),
.SAXIGP5WREADY (pl_to_ps_axi_hp3_fpd_wready),
.SAXIGP5BID (pl_to_ps_axi_hp3_fpd_bid),
.SAXIGP5BRESP (pl_to_ps_axi_hp3_fpd_bresp),
.SAXIGP5BVALID (pl_to_ps_axi_hp3_fpd_bvalid),
.SAXIGP5BREADY (pl_to_ps_axi_hp3_fpd_bready),
.SAXIGP5ARID (pl_to_ps_axi_hp3_fpd_arid),
.SAXIGP5ARADDR (pl_to_ps_axi_hp3_fpd_araddr),
.SAXIGP5ARLEN (pl_to_ps_axi_hp3_fpd_arlen),
.SAXIGP5ARSIZE (pl_to_ps_axi_hp3_fpd_arsize),
.SAXIGP5ARBURST (pl_to_ps_axi_hp3_fpd_arburst),
.SAXIGP5ARLOCK (pl_to_ps_axi_hp3_fpd_arlock),
.SAXIGP5ARCACHE (pl_to_ps_axi_hp3_fpd_arcache),
.SAXIGP5ARPROT (pl_to_ps_axi_hp3_fpd_arprot),
.SAXIGP5ARVALID (pl_to_ps_axi_hp3_fpd_arvalid),
.SAXIGP5ARREADY (pl_to_ps_axi_hp3_fpd_arready),
.SAXIGP5RID (pl_to_ps_axi_hp3_fpd_rid),
.SAXIGP5RDATA (pl_to_ps_axi_hp3_fpd_rdata),
.SAXIGP5RRESP (pl_to_ps_axi_hp3_fpd_rresp),
.SAXIGP5RLAST (pl_to_ps_axi_hp3_fpd_rlast),
.SAXIGP5RVALID (pl_to_ps_axi_hp3_fpd_rvalid),
.SAXIGP5RREADY (pl_to_ps_axi_hp3_fpd_rready),
.SAXIGP5AWQOS (pl_to_ps_axi_hp3_fpd_awqos),
.SAXIGP5ARQOS (pl_to_ps_axi_hp3_fpd_arqos),
.SAXIGP5RCOUNT (pl_to_ps_axi_hp3_fpd_rcount),
.SAXIGP5WCOUNT (pl_to_ps_axi_hp3_fpd_wcount),
.SAXIGP5RACOUNT (pl_to_ps_axi_hp3_fpd_racount),
.SAXIGP5WACOUNT (pl_to_ps_axi_hp3_fpd_wacount),
.SAXIGP6RCLK (clk_pl_to_ps_axi_lpd_read),
.SAXIGP6WCLK (clk_pl_to_ps_axi_lpd_write),
.SAXIGP6ARUSER (pl_to_ps_axi_lpd_aruser),
.SAXIGP6AWUSER (pl_to_ps_axi_lpd_awuser),
.SAXIGP6AWID (pl_to_ps_axi_lpd_awid),
.SAXIGP6AWADDR (pl_to_ps_axi_lpd_awaddr),
.SAXIGP6AWLEN (pl_to_ps_axi_lpd_awlen),
.SAXIGP6AWSIZE (pl_to_ps_axi_lpd_awsize),
.SAXIGP6AWBURST (pl_to_ps_axi_lpd_awburst),
.SAXIGP6AWLOCK (pl_to_ps_axi_lpd_awlock),
.SAXIGP6AWCACHE (pl_to_ps_axi_lpd_awcache),
.SAXIGP6AWPROT (pl_to_ps_axi_lpd_awprot),
.SAXIGP6AWVALID (pl_to_ps_axi_lpd_awvalid),
.SAXIGP6AWREADY (pl_to_ps_axi_lpd_awready),
.SAXIGP6WDATA (pl_to_ps_axi_lpd_wdata),
.SAXIGP6WSTRB (pl_to_ps_axi_lpd_wstrb),
.SAXIGP6WLAST (pl_to_ps_axi_lpd_wlast),
.SAXIGP6WVALID (pl_to_ps_axi_lpd_wvalid),
.SAXIGP6WREADY (pl_to_ps_axi_lpd_wready),
.SAXIGP6BID (pl_to_ps_axi_lpd_bid),
.SAXIGP6BRESP (pl_to_ps_axi_lpd_bresp),
.SAXIGP6BVALID (pl_to_ps_axi_lpd_bvalid),
.SAXIGP6BREADY (pl_to_ps_axi_lpd_bready),
.SAXIGP6ARID (pl_to_ps_axi_lpd_arid),
.SAXIGP6ARADDR (pl_to_ps_axi_lpd_araddr),
.SAXIGP6ARLEN (pl_to_ps_axi_lpd_arlen),
.SAXIGP6ARSIZE (pl_to_ps_axi_lpd_arsize),
.SAXIGP6ARBURST (pl_to_ps_axi_lpd_arburst),
.SAXIGP6ARLOCK (pl_to_ps_axi_lpd_arlock),
.SAXIGP6ARCACHE (pl_to_ps_axi_lpd_arcache),
.SAXIGP6ARPROT (pl_to_ps_axi_lpd_arprot),
.SAXIGP6ARVALID (pl_to_ps_axi_lpd_arvalid),
.SAXIGP6ARREADY (pl_to_ps_axi_lpd_arready),
.SAXIGP6RID (pl_to_ps_axi_lpd_rid),
.SAXIGP6RDATA (pl_to_ps_axi_lpd_rdata),
.SAXIGP6RRESP (pl_to_ps_axi_lpd_rresp),
.SAXIGP6RLAST (pl_to_ps_axi_lpd_rlast),
.SAXIGP6RVALID (pl_to_ps_axi_lpd_rvalid),
.SAXIGP6RREADY (pl_to_ps_axi_lpd_rready),
.SAXIGP6AWQOS (pl_to_ps_axi_lpd_awqos),
.SAXIGP6ARQOS (pl_to_ps_axi_lpd_arqos),
.SAXIGP6RCOUNT (pl_to_ps_axi_lpd_rcount),
.SAXIGP6WCOUNT (pl_to_ps_axi_lpd_wcount),
.SAXIGP6RACOUNT (pl_to_ps_axi_lpd_racount),
.SAXIGP6WACOUNT (pl_to_ps_axi_lpd_wacount),
.SAXIACPACLK (clk_pl_to_ps_consumer_acp_fpd),
.SAXIACPAWADDR (pl_to_ps_axi_acp_fpd_awaddr),
.SAXIACPAWID (pl_to_ps_axi_acp_fpd_awid),
.SAXIACPAWLEN (pl_to_ps_axi_acp_fpd_awlen),
.SAXIACPAWSIZE (pl_to_ps_axi_acp_fpd_awsize),
.SAXIACPAWBURST (pl_to_ps_axi_acp_fpd_awburst),
.SAXIACPAWLOCK (pl_to_ps_axi_acp_fpd_awlock),
.SAXIACPAWCACHE (pl_to_ps_axi_acp_fpd_awcache),
.SAXIACPAWPROT (pl_to_ps_axi_acp_fpd_awprot),
.SAXIACPAWVALID (pl_to_ps_axi_acp_fpd_awvalid),
.SAXIACPAWREADY (pl_to_ps_axi_acp_fpd_awready),
.SAXIACPAWUSER (pl_to_ps_axi_acp_fpd_awuser),
.SAXIACPAWQOS (pl_to_ps_axi_acp_fpd_awqos),
.SAXIACPWLAST (pl_to_ps_axi_acp_fpd_wlast),
.SAXIACPWDATA (pl_to_ps_axi_acp_fpd_wdata),
.SAXIACPWSTRB (pl_to_ps_axi_acp_fpd_wstrb),
.SAXIACPWVALID (pl_to_ps_axi_acp_fpd_wvalid),
.SAXIACPWREADY (pl_to_ps_axi_acp_fpd_wready),
.SAXIACPBRESP (pl_to_ps_axi_acp_fpd_bresp),
.SAXIACPBID (pl_to_ps_axi_acp_fpd_bid),
.SAXIACPBVALID (pl_to_ps_axi_acp_fpd_bvalid),
.SAXIACPBREADY (pl_to_ps_axi_acp_fpd_bready),
.SAXIACPARADDR (pl_to_ps_axi_acp_fpd_araddr),
.SAXIACPARID (pl_to_ps_axi_acp_fpd_arid),
.SAXIACPARLEN (pl_to_ps_axi_acp_fpd_arlen),
.SAXIACPARSIZE (pl_to_ps_axi_acp_fpd_arsize),
.SAXIACPARBURST (pl_to_ps_axi_acp_fpd_arburst),
.SAXIACPARLOCK (pl_to_ps_axi_acp_fpd_arlock),
.SAXIACPARCACHE (pl_to_ps_axi_acp_fpd_arcache),
.SAXIACPARPROT (pl_to_ps_axi_acp_fpd_arprot),
.SAXIACPARVALID (pl_to_ps_axi_acp_fpd_arvalid),
.SAXIACPARREADY (pl_to_ps_axi_acp_fpd_arready),
.SAXIACPARUSER (pl_to_ps_axi_acp_fpd_aruser),
.SAXIACPARQOS (pl_to_ps_axi_acp_fpd_arqos),
.SAXIACPRID (pl_to_ps_axi_acp_fpd_rid),
.SAXIACPRLAST (pl_to_ps_axi_acp_fpd_rlast),
.SAXIACPRDATA (pl_to_ps_axi_acp_fpd_rdata),
.SAXIACPRRESP (pl_to_ps_axi_acp_fpd_rresp),
.SAXIACPRVALID (pl_to_ps_axi_acp_fpd_rvalid),
.SAXIACPRREADY (pl_to_ps_axi_acp_fpd_rready),
.PLACECLK (pl_to_ps_axi_ace_fpd_aclk),
.SACEFPDAWVALID (pl_to_ps_axi_ace_fpd_awvalid),
.SACEFPDAWREADY (pl_to_ps_axi_ace_fpd_awready),
.SACEFPDAWID (pl_to_ps_axi_ace_fpd_awid),
.SACEFPDAWADDR (pl_to_ps_axi_ace_fpd_awaddr),
.SACEFPDAWREGION (pl_to_ps_axi_ace_fpd_awregion),
.SACEFPDAWLEN (pl_to_ps_axi_ace_fpd_awlen),
.SACEFPDAWSIZE (pl_to_ps_axi_ace_fpd_awsize),
.SACEFPDAWBURST (pl_to_ps_axi_ace_fpd_awburst),
.SACEFPDAWLOCK (pl_to_ps_axi_ace_fpd_awlock),
.SACEFPDAWCACHE (pl_to_ps_axi_ace_fpd_awcache),
.SACEFPDAWPROT (pl_to_ps_axi_ace_fpd_awprot),
.SACEFPDAWDOMAIN (pl_to_ps_axi_ace_fpd_awdomain),
.SACEFPDAWSNOOP (pl_to_ps_axi_ace_fpd_awsnoop),
.SACEFPDAWBAR (pl_to_ps_axi_ace_fpd_awbar),
.SACEFPDAWQOS (pl_to_ps_axi_ace_fpd_awqos),
.SACEFPDAWUSER (pl_to_ps_axi_ace_fpd_awuser),
.SACEFPDWVALID (pl_to_ps_axi_ace_fpd_wvalid),
.SACEFPDWREADY (pl_to_ps_axi_ace_fpd_wready),
.SACEFPDWDATA (pl_to_ps_axi_ace_fpd_wdata),
.SACEFPDWSTRB (pl_to_ps_axi_ace_fpd_wstrb),
.SACEFPDWLAST (pl_to_ps_axi_ace_fpd_wlast),
.SACEFPDWUSER (pl_to_ps_axi_ace_fpd_wuser),
.SACEFPDBVALID (pl_to_ps_axi_ace_fpd_bvalid),
.SACEFPDBREADY (pl_to_ps_axi_ace_fpd_bready),
.SACEFPDBID (pl_to_ps_axi_ace_fpd_bid),
.SACEFPDBRESP (pl_to_ps_axi_ace_fpd_bresp),
.SACEFPDBUSER (pl_to_ps_axi_ace_fpd_buser),
.SACEFPDARVALID (pl_to_ps_axi_ace_fpd_arvalid),
.SACEFPDARREADY (pl_to_ps_axi_ace_fpd_arready),
.SACEFPDARID (pl_to_ps_axi_ace_fpd_arid),
.SACEFPDARADDR (pl_to_ps_axi_ace_fpd_araddr),
.SACEFPDARREGION (pl_to_ps_axi_ace_fpd_arregion),
.SACEFPDARLEN (pl_to_ps_axi_ace_fpd_arlen),
.SACEFPDARSIZE (pl_to_ps_axi_ace_fpd_arsize),
.SACEFPDARBURST (pl_to_ps_axi_ace_fpd_arburst),
.SACEFPDARLOCK (pl_to_ps_axi_ace_fpd_arlock),
.SACEFPDARCACHE (pl_to_ps_axi_ace_fpd_arcache),
.SACEFPDARPROT (pl_to_ps_axi_ace_fpd_arprot),
.SACEFPDARDOMAIN (pl_to_ps_axi_ace_fpd_ardomain),
.SACEFPDARSNOOP (pl_to_ps_axi_ace_fpd_arsnoop),
.SACEFPDARBAR (pl_to_ps_axi_ace_fpd_arbar),
.SACEFPDARQOS (pl_to_ps_axi_ace_fpd_arqos),
.SACEFPDARUSER (pl_to_ps_axi_ace_fpd_aruser),
.SACEFPDRVALID (pl_to_ps_axi_ace_fpd_rvalid),
.SACEFPDRREADY (pl_to_ps_axi_ace_fpd_rready),
.SACEFPDRID (pl_to_ps_axi_ace_fpd_rid),
.SACEFPDRDATA (pl_to_ps_axi_ace_fpd_rdata),
.SACEFPDRRESP (pl_to_ps_axi_ace_fpd_rresp),
.SACEFPDRLAST (pl_to_ps_axi_ace_fpd_rlast),
.SACEFPDRUSER (pl_to_ps_axi_ace_fpd_ruser),
.SACEFPDACVALID (pl_to_ps_axi_ace_fpd_acvalid),
.SACEFPDACREADY (pl_to_ps_axi_ace_fpd_acready),
.SACEFPDACADDR (pl_to_ps_axi_ace_fpd_acaddr),
.SACEFPDACSNOOP (pl_to_ps_axi_ace_fpd_acsnoop),
.SACEFPDACPROT (pl_to_ps_axi_ace_fpd_acprot),
.SACEFPDCRVALID (pl_to_ps_axi_ace_fpd_crvalid),
.SACEFPDCRREADY (pl_to_ps_axi_ace_fpd_crready),
.SACEFPDCRRESP (pl_to_ps_axi_ace_fpd_crresp),
.SACEFPDCDVALID (pl_to_ps_axi_ace_fpd_cdvalid),
.SACEFPDCDREADY (pl_to_ps_axi_ace_fpd_cdready),
.SACEFPDCDDATA (pl_to_ps_axi_ace_fpd_cddata),
.SACEFPDCDLAST (pl_to_ps_axi_ace_fpd_cdlast),
.SACEFPDWACK (pl_to_ps_axi_ace_fpd_wack),
.SACEFPDRACK (pl_to_ps_axi_ace_fpd_rack),
.EMIOCAN0PHYTX (emio_can0_phy_tx),
.EMIOCAN0PHYRX (emio_can0_phy_rx),
.EMIOCAN1PHYTX (emio_can1_phy_tx),
.EMIOCAN1PHYRX (emio_can1_phy_rx),
.EMIOENET0GMIIRXCLK (clk_pl_to_ps_emio_enet0_gmii_rx),
.EMIOENET0SPEEDMODE (emio_enet0_speed_mode),
.EMIOENET0GMIICRS (emio_enet0_gmii_crs),
.EMIOENET0GMIICOL (emio_enet0_gmii_col),
.EMIOENET0GMIIRXD (emio_enet0_gmii_rxd),
.EMIOENET0GMIIRXER (emio_enet0_gmii_rx_er),
.EMIOENET0GMIIRXDV (emio_enet0_gmii_rx_dv),
.EMIOENET0GMIITXCLK (clk_pl_to_ps_emio_enet0_gmii_tx),
.EMIOENET0GMIITXD (emio_enet0_gmii_txd),
.EMIOENET0GMIITXEN (emio_enet0_gmii_tx_en),
.EMIOENET0GMIITXER (emio_enet0_gmii_tx_er),
.EMIOENET0MDIOMDC (emio_enet0_mdio_mdc),
.EMIOENET0MDIOI (emio_enet0_mdio_i),
.EMIOENET0MDIOO (emio_enet0_mdio_o),
.EMIOENET0MDIOTN (emio_enet0_mdio_t_n),
.EMIOENET1GMIIRXCLK (clk_pl_to_ps_emio_enet1_gmii_rx),
.EMIOENET1SPEEDMODE (emio_enet1_speed_mode),
.EMIOENET1GMIICRS (emio_enet1_gmii_crs),
.EMIOENET1GMIICOL (emio_enet1_gmii_col),
.EMIOENET1GMIIRXD (emio_enet1_gmii_rxd),
.EMIOENET1GMIIRXER (emio_enet1_gmii_rx_er),
.EMIOENET1GMIIRXDV (emio_enet1_gmii_rx_dv),
.EMIOENET1GMIITXCLK (clk_pl_to_ps_emio_enet1_gmii_tx),
.EMIOENET1GMIITXD (emio_enet1_gmii_txd),
.EMIOENET1GMIITXEN (emio_enet1_gmii_tx_en),
.EMIOENET1GMIITXER (emio_enet1_gmii_tx_er),
.EMIOENET1MDIOMDC (emio_enet1_mdio_mdc),
.EMIOENET1MDIOI (emio_enet1_mdio_i),
.EMIOENET1MDIOO (emio_enet1_mdio_o),
.EMIOENET1MDIOTN (emio_enet1_mdio_t_n),
.EMIOENET2GMIIRXCLK (clk_pl_to_ps_emio_enet2_gmii_rx),
.EMIOENET2SPEEDMODE (emio_enet2_speed_mode),
.EMIOENET2GMIICRS (emio_enet2_gmii_crs),
.EMIOENET2GMIICOL (emio_enet2_gmii_col),
.EMIOENET2GMIIRXD (emio_enet2_gmii_rxd),
.EMIOENET2GMIIRXER (emio_enet2_gmii_rx_er),
.EMIOENET2GMIIRXDV (emio_enet2_gmii_rx_dv),
.EMIOENET2GMIITXCLK (clk_pl_to_ps_emio_enet2_gmii_tx),
.EMIOENET2GMIITXD (emio_enet2_gmii_txd),
.EMIOENET2GMIITXEN (emio_enet2_gmii_tx_en),
.EMIOENET2GMIITXER (emio_enet2_gmii_tx_er),
.EMIOENET2MDIOMDC (emio_enet2_mdio_mdc),
.EMIOENET2MDIOI (emio_enet2_mdio_i),
.EMIOENET2MDIOO (emio_enet2_mdio_o),
.EMIOENET2MDIOTN (emio_enet2_mdio_t_n),
.EMIOENET3GMIIRXCLK (clk_pl_to_ps_emio_enet3_gmii_rx),
.EMIOENET3SPEEDMODE (emio_enet3_speed_mode),
.EMIOENET3GMIICRS (emio_enet3_gmii_crs),
.EMIOENET3GMIICOL (emio_enet3_gmii_col),
.EMIOENET3GMIIRXD (emio_enet3_gmii_rxd),
.EMIOENET3GMIIRXER (emio_enet3_gmii_rx_er),
.EMIOENET3GMIIRXDV (emio_enet3_gmii_rx_dv),
.EMIOENET3GMIITXCLK (clk_pl_to_ps_emio_enet3_gmii_tx),
.EMIOENET3GMIITXD (emio_enet3_gmii_txd),
.EMIOENET3GMIITXEN (emio_enet3_gmii_tx_en),
.EMIOENET3GMIITXER (emio_enet3_gmii_tx_er),
.EMIOENET3MDIOMDC (emio_enet3_mdio_mdc),
.EMIOENET3MDIOI (emio_enet3_mdio_i),
.EMIOENET3MDIOO (emio_enet3_mdio_o),
.EMIOENET3MDIOTN (emio_enet3_mdio_t_n),
.EMIOENET0TXRDATARDY (emio_enet0_tx_r_data_rdy),
.EMIOENET0TXRRD (emio_enet0_tx_r_rd),
.EMIOENET0TXRVALID (emio_enet0_tx_r_valid),
.EMIOENET0TXRDATA (emio_enet0_tx_r_data),
.EMIOENET0TXRSOP (emio_enet0_tx_r_sop),
.EMIOENET0TXREOP (emio_enet0_tx_r_eop),
.EMIOENET0TXRERR (emio_enet0_tx_r_err),
.EMIOENET0TXRUNDERFLOW (emio_enet0_tx_r_underflow),
.EMIOENET0TXRFLUSHED (emio_enet0_tx_r_flushed),
.EMIOENET0TXRCONTROL (emio_enet0_tx_r_control),
.EMIOENET0DMATXENDTOG (emio_enet0_dma_tx_end_tog),
.EMIOENET0DMATXSTATUSTOG (emio_enet0_dma_tx_status_tog),
.EMIOENET0TXRSTATUS (emio_enet0_tx_r_status),
.EMIOENET0RXWWR (emio_enet0_rx_w_wr),
.EMIOENET0RXWDATA (emio_enet0_rx_w_data),
.EMIOENET0RXWSOP (emio_enet0_rx_w_sop),
.EMIOENET0RXWEOP (emio_enet0_rx_w_eop),
.EMIOENET0RXWSTATUS (emio_enet0_rx_w_status),
.EMIOENET0RXWERR (emio_enet0_rx_w_err),
.EMIOENET0RXWOVERFLOW (emio_enet0_rx_w_overflow),
.FMIOGEM0SIGNALDETECT (emio_enet0_signal_detect),
.EMIOENET0RXWFLUSH (emio_enet0_rx_w_flush),
.EMIOGEM0TXRFIXEDLAT (emio_enet0_tx_r_fixed_lat),
.FMIOGEM0FIFOTXCLKFROMPL (clk_pl_to_ps_fmio_gem0_fifo_tx),
.FMIOGEM0FIFORXCLKFROMPL (clk_pl_to_ps_fmio_gem0_fifo_rx),
.FMIOGEM0FIFOTXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem0_fifo_tx),
.FMIOGEM0FIFORXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem0_fifo_rx),
.EMIOENET1TXRDATARDY (emio_enet1_tx_r_data_rdy),
.EMIOENET1TXRRD (emio_enet1_tx_r_rd),
.EMIOENET1TXRVALID (emio_enet1_tx_r_valid),
.EMIOENET1TXRDATA (emio_enet1_tx_r_data),
.EMIOENET1TXRSOP (emio_enet1_tx_r_sop),
.EMIOENET1TXREOP (emio_enet1_tx_r_eop),
.EMIOENET1TXRERR (emio_enet1_tx_r_err),
.EMIOENET1TXRUNDERFLOW (emio_enet1_tx_r_underflow),
.EMIOENET1TXRFLUSHED (emio_enet1_tx_r_flushed),
.EMIOENET1TXRCONTROL (emio_enet1_tx_r_control),
.EMIOENET1DMATXENDTOG (emio_enet1_dma_tx_end_tog),
.EMIOENET1DMATXSTATUSTOG (emio_enet1_dma_tx_status_tog),
.EMIOENET1TXRSTATUS (emio_enet1_tx_r_status),
.EMIOENET1RXWWR (emio_enet1_rx_w_wr),
.EMIOENET1RXWDATA (emio_enet1_rx_w_data),
.EMIOENET1RXWSOP (emio_enet1_rx_w_sop),
.EMIOENET1RXWEOP (emio_enet1_rx_w_eop),
.EMIOENET1RXWSTATUS (emio_enet1_rx_w_status),
.EMIOENET1RXWERR (emio_enet1_rx_w_err),
.EMIOENET1RXWOVERFLOW (emio_enet1_rx_w_overflow),
.FMIOGEM1SIGNALDETECT (emio_enet1_signal_detect),
.EMIOENET1RXWFLUSH (emio_enet1_rx_w_flush),
.EMIOGEM1TXRFIXEDLAT (emio_enet1_tx_r_fixed_lat),
.FMIOGEM1FIFOTXCLKFROMPL (clk_pl_to_ps_fmio_gem1_fifo_tx),
.FMIOGEM1FIFORXCLKFROMPL (clk_pl_to_ps_fmio_gem1_fifo_rx),
.FMIOGEM1FIFOTXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem1_fifo_tx),
.FMIOGEM1FIFORXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem1_fifo_rx),
.EMIOENET2TXRDATARDY (emio_enet2_tx_r_data_rdy),
.EMIOENET2TXRRD (emio_enet2_tx_r_rd),
.EMIOENET2TXRVALID (emio_enet2_tx_r_valid),
.EMIOENET2TXRDATA (emio_enet2_tx_r_data),
.EMIOENET2TXRSOP (emio_enet2_tx_r_sop),
.EMIOENET2TXREOP (emio_enet2_tx_r_eop),
.EMIOENET2TXRERR (emio_enet2_tx_r_err),
.EMIOENET2TXRUNDERFLOW (emio_enet2_tx_r_underflow),
.EMIOENET2TXRFLUSHED (emio_enet2_tx_r_flushed),
.EMIOENET2TXRCONTROL (emio_enet2_tx_r_control),
.EMIOENET2DMATXENDTOG (emio_enet2_dma_tx_end_tog),
.EMIOENET2DMATXSTATUSTOG (emio_enet2_dma_tx_status_tog),
.EMIOENET2TXRSTATUS (emio_enet2_tx_r_status),
.EMIOENET2RXWWR (emio_enet2_rx_w_wr),
.EMIOENET2RXWDATA (emio_enet2_rx_w_data),
.EMIOENET2RXWSOP (emio_enet2_rx_w_sop),
.EMIOENET2RXWEOP (emio_enet2_rx_w_eop),
.EMIOENET2RXWSTATUS (emio_enet2_rx_w_status),
.EMIOENET2RXWERR (emio_enet2_rx_w_err),
.EMIOENET2RXWOVERFLOW (emio_enet2_rx_w_overflow),
.FMIOGEM2SIGNALDETECT (emio_enet2_signal_detect),
.EMIOENET2RXWFLUSH (emio_enet2_rx_w_flush),
.EMIOGEM2TXRFIXEDLAT (emio_enet2_tx_r_fixed_lat),
.FMIOGEM2FIFOTXCLKFROMPL (clk_pl_to_ps_fmio_gem2_fifo_tx),
.FMIOGEM2FIFORXCLKFROMPL (clk_pl_to_ps_fmio_gem2_fifo_rx),
.FMIOGEM2FIFOTXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem2_fifo_tx),
.FMIOGEM2FIFORXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem2_fifo_rx),
.EMIOENET3TXRDATARDY (emio_enet3_tx_r_data_rdy),
.EMIOENET3TXRRD (emio_enet3_tx_r_rd),
.EMIOENET3TXRVALID (emio_enet3_tx_r_valid),
.EMIOENET3TXRDATA (emio_enet3_tx_r_data),
.EMIOENET3TXRSOP (emio_enet3_tx_r_sop),
.EMIOENET3TXREOP (emio_enet3_tx_r_eop),
.EMIOENET3TXRERR (emio_enet3_tx_r_err),
.EMIOENET3TXRUNDERFLOW (emio_enet3_tx_r_underflow),
.EMIOENET3TXRFLUSHED (emio_enet3_tx_r_flushed),
.EMIOENET3TXRCONTROL (emio_enet3_tx_r_control),
.EMIOENET3DMATXENDTOG (emio_enet3_dma_tx_end_tog),
.EMIOENET3DMATXSTATUSTOG (emio_enet3_dma_tx_status_tog),
.EMIOENET3TXRSTATUS (emio_enet3_tx_r_status),
.EMIOENET3RXWWR (emio_enet3_rx_w_wr),
.EMIOENET3RXWDATA (emio_enet3_rx_w_data),
.EMIOENET3RXWSOP (emio_enet3_rx_w_sop),
.EMIOENET3RXWEOP (emio_enet3_rx_w_eop),
.EMIOENET3RXWSTATUS (emio_enet3_rx_w_status),
.EMIOENET3RXWERR (emio_enet3_rx_w_err),
.EMIOENET3RXWOVERFLOW (emio_enet3_rx_w_overflow),
.FMIOGEM3SIGNALDETECT (emio_enet3_signal_detect),
.EMIOENET3RXWFLUSH (emio_enet3_rx_w_flush),
.EMIOGEM3TXRFIXEDLAT (emio_enet3_tx_r_fixed_lat),
.FMIOGEM3FIFOTXCLKFROMPL (clk_pl_to_ps_fmio_gem3_fifo_tx),
.FMIOGEM3FIFORXCLKFROMPL (clk_pl_to_ps_fmio_gem3_fifo_rx),
.FMIOGEM3FIFOTXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem3_fifo_tx),
.FMIOGEM3FIFORXCLKTOPLBUFG (clk_ps_to_pl_fmio_gem3_fifo_rx),
.EMIOGEM0TXSOF (emio_enet0_tx_sof),
.EMIOGEM0SYNCFRAMETX (emio_enet0_sync_frame_tx),
.EMIOGEM0DELAYREQTX (emio_enet0_delay_req_tx),
.EMIOGEM0PDELAYREQTX (emio_enet0_pdelay_req_tx),
.EMIOGEM0PDELAYRESPTX (emio_enet0_pdelay_resp_tx),
.EMIOGEM0RXSOF (emio_enet0_rx_sof),
.EMIOGEM0SYNCFRAMERX (emio_enet0_sync_frame_rx),
.EMIOGEM0DELAYREQRX (emio_enet0_delay_req_rx),
.EMIOGEM0PDELAYREQRX (emio_enet0_pdelay_req_rx),
.EMIOGEM0PDELAYRESPRX (emio_enet0_pdelay_resp_rx),
.EMIOGEM0TSUINCCTRL (emio_enet0_tsu_inc_ctrl),
.EMIOGEM0TSUTIMERCMPVAL (emio_enet0_tsu_timer_cmp_val),
.EMIOGEM1TXSOF (emio_enet1_tx_sof),
.EMIOGEM1SYNCFRAMETX (emio_enet1_sync_frame_tx),
.EMIOGEM1DELAYREQTX (emio_enet1_delay_req_tx),
.EMIOGEM1PDELAYREQTX (emio_enet1_pdelay_req_tx),
.EMIOGEM1PDELAYRESPTX (emio_enet1_pdelay_resp_tx),
.EMIOGEM1RXSOF (emio_enet1_rx_sof),
.EMIOGEM1SYNCFRAMERX (emio_enet1_sync_frame_rx),
.EMIOGEM1DELAYREQRX (emio_enet1_delay_req_rx),
.EMIOGEM1PDELAYREQRX (emio_enet1_pdelay_req_rx),
.EMIOGEM1PDELAYRESPRX (emio_enet1_pdelay_resp_rx),
.EMIOGEM1TSUINCCTRL (emio_enet1_tsu_inc_ctrl),
.EMIOGEM1TSUTIMERCMPVAL (emio_enet1_tsu_timer_cmp_val),
.EMIOGEM2TXSOF (emio_enet2_tx_sof),
.EMIOGEM2SYNCFRAMETX (emio_enet2_sync_frame_tx),
.EMIOGEM2DELAYREQTX (emio_enet2_delay_req_tx),
.EMIOGEM2PDELAYREQTX (emio_enet2_pdelay_req_tx),
.EMIOGEM2PDELAYRESPTX (emio_enet2_pdelay_resp_tx),
.EMIOGEM2RXSOF (emio_enet2_rx_sof),
.EMIOGEM2SYNCFRAMERX (emio_enet2_sync_frame_rx),
.EMIOGEM2DELAYREQRX (emio_enet2_delay_req_rx),
.EMIOGEM2PDELAYREQRX (emio_enet2_pdelay_req_rx),
.EMIOGEM2PDELAYRESPRX (emio_enet2_pdelay_resp_rx),
.EMIOGEM2TSUINCCTRL (emio_enet2_tsu_inc_ctrl),
.EMIOGEM2TSUTIMERCMPVAL (emio_enet2_tsu_timer_cmp_val),
.EMIOGEM3TXSOF (emio_enet3_tx_sof),
.EMIOGEM3SYNCFRAMETX (emio_enet3_sync_frame_tx),
.EMIOGEM3DELAYREQTX (emio_enet3_delay_req_tx),
.EMIOGEM3PDELAYREQTX (emio_enet3_pdelay_req_tx),
.EMIOGEM3PDELAYRESPTX (emio_enet3_pdelay_resp_tx),
.EMIOGEM3RXSOF (emio_enet3_rx_sof),
.EMIOGEM3SYNCFRAMERX (emio_enet3_sync_frame_rx),
.EMIOGEM3DELAYREQRX (emio_enet3_delay_req_rx),
.EMIOGEM3PDELAYREQRX (emio_enet3_pdelay_req_rx),
.EMIOGEM3PDELAYRESPRX (emio_enet3_pdelay_resp_rx),
.EMIOGEM3TSUINCCTRL (emio_enet3_tsu_inc_ctrl),
.EMIOGEM3TSUTIMERCMPVAL (emio_enet3_tsu_timer_cmp_val),
.FMIOGEMTSUCLKFROMPL (clk_pl_to_ps_fmio_gem_tsu),
.FMIOGEMTSUCLKTOPLBUFG (clk_ps_to_pl_gem_tsu_clk),
.EMIOENETTSUCLK (clk_pl_to_ps_emio_enet_tsu),
.EMIOENET0GEMTSUTIMERCNT (emio_enet0_enet_tsu_timer_cnt),
.EMIOENET0EXTINTIN (emio_enet0_ext_int_in),
.EMIOENET1EXTINTIN (emio_enet1_ext_int_in),
.EMIOENET2EXTINTIN (emio_enet2_ext_int_in),
.EMIOENET3EXTINTIN (emio_enet3_ext_int_in),
.EMIOENET0DMABUSWIDTH (emio_enet0_dma_bus_width),
.EMIOENET1DMABUSWIDTH (emio_enet1_dma_bus_width),
.EMIOENET2DMABUSWIDTH (emio_enet2_dma_bus_width),
.EMIOENET3DMABUSWIDTH (emio_enet3_dma_bus_width),
.EMIOGPIOI (emio_gpio_i),
.EMIOGPIOO (emio_gpio_o),
.EMIOGPIOTN (emio_gpio_t_n),
.EMIOI2C0SCLI (emio_i2c0_scl_i),
.EMIOI2C0SCLO (emio_i2c0_scl_o),
.EMIOI2C0SCLTN (emio_i2c0_scl_tri),
.EMIOI2C0SDAI (emio_i2c0_sda_i),
.EMIOI2C0SDAO (emio_i2c0_sda_o),
.EMIOI2C0SDATN (emio_i2c0_sda_t_n),
.EMIOI2C1SCLI (emio_i2c1_scl_i),
.EMIOI2C1SCLO (emio_i2c1_scl_o),
.EMIOI2C1SCLTN (emio_i2c1_scl_tri),
.EMIOI2C1SDAI (emio_i2c1_sda_i),
.EMIOI2C1SDAO (emio_i2c1_sda_o),
.EMIOI2C1SDATN (emio_i2c1_sda_t_n),
.EMIOUART0TX (emio_uart0_txd),
.EMIOUART0RX (emio_uart0_rxd),
.EMIOUART0CTSN (emio_uart0_ctsn),
.EMIOUART0RTSN (emio_uart0_rtsn),
.EMIOUART0DSRN (emio_uart0_dsrn),
.EMIOUART0DCDN (emio_uart0_dcdn),
.EMIOUART0RIN (emio_uart0_rin),
.EMIOUART0DTRN (emio_uart0_dtrn),
.EMIOUART1TX (emio_uart1_txd),
.EMIOUART1RX (emio_uart1_rxd),
.EMIOUART1CTSN (emio_uart1_ctsn),
.EMIOUART1RTSN (emio_uart1_rtsn),
.EMIOUART1DSRN (emio_uart1_dsrn),
.EMIOUART1DCDN (emio_uart1_dcdn),
.EMIOUART1RIN (emio_uart1_rin),
.EMIOUART1DTRN (emio_uart1_dtrn),
.EMIOSDIO0CLKOUT (clk_ps_to_pl_emio_sdio0),
.EMIOSDIO0FBCLKIN (clk_pl_to_ps_emio_sdio0),
.EMIOSDIO0CMDOUT (emio_sdio0_cmdout),
.EMIOSDIO0CMDIN (emio_sdio0_cmdin),
.EMIOSDIO0CMDENA (emio_sdio0_cmdena_n),
.EMIOSDIO0DATAIN (emio_sdio0_datain),
.EMIOSDIO0DATAOUT (emio_sdio0_dataout),
.EMIOSDIO0DATAENA (emio_sdio0_dataena_n),
.EMIOSDIO0CDN (emio_sdio0_cd_n),
.EMIOSDIO0WP (emio_sdio0_wp),
.EMIOSDIO0LEDCONTROL (emio_sdio0_ledcontrol),
.EMIOSDIO0BUSPOWER (emio_sdio0_buspower),
.EMIOSDIO0BUSVOLT (emio_sdio0_bus_volt),
.EMIOSDIO1CLKOUT (clk_ps_to_pl_emio_sdio1),
.EMIOSDIO1FBCLKIN (clk_pl_to_ps_emio_sdio1),
.EMIOSDIO1CMDOUT (emio_sdio1_cmdout),
.EMIOSDIO1CMDIN (emio_sdio1_cmdin),
.EMIOSDIO1CMDENA (emio_sdio1_cmdena_n),
.EMIOSDIO1DATAIN (emio_sdio1_datain),
.EMIOSDIO1DATAOUT (emio_sdio1_dataout),
.EMIOSDIO1DATAENA (emio_sdio1_dataena_n),
.EMIOSDIO1CDN (emio_sdio1_cd_n),
.EMIOSDIO1WP (emio_sdio1_wp),
.EMIOSDIO1LEDCONTROL (emio_sdio1_ledcontrol),
.EMIOSDIO1BUSPOWER (emio_sdio1_buspower),
.EMIOSDIO1BUSVOLT (emio_sdio1_bus_volt),
.EMIOSPI0SCLKI (emio_spi0_sclk_i),
.EMIOSPI0SCLKO (emio_spi0_sclk_o),
.EMIOSPI0SCLKTN (emio_spi0_sclk_t_n),
.EMIOSPI0MI (emio_spi0_m_i),
.EMIOSPI0MO (emio_spi0_m_o),
.EMIOSPI0MOTN (emio_spi0_mo_t_n),
.EMIOSPI0SI (emio_spi0_s_i),
.EMIOSPI0SO (emio_spi0_s_o),
.EMIOSPI0STN (emio_spi0_so_t_n),
.EMIOSPI0SSIN (emio_spi0_ss_i_n),
.EMIOSPI0SSON ({emio_spi0_ss2_o_n,emio_spi0_ss1_o_n,emio_spi0_ss_o_n}),
.EMIOSPI0SSNTN (emio_spi0_ss_n_t_n),
.EMIOSPI1SCLKI (emio_spi1_sclk_i),
.EMIOSPI1SCLKO (emio_spi1_sclk_o),
.EMIOSPI1SCLKTN (emio_spi1_sclk_t_n),
.EMIOSPI1MI (emio_spi1_m_i),
.EMIOSPI1MO (emio_spi1_m_o),
.EMIOSPI1MOTN (emio_spi1_mo_t_n),
.EMIOSPI1SI (emio_spi1_s_i),
.EMIOSPI1SO (emio_spi1_s_o),
.EMIOSPI1STN (emio_spi1_so_tri),
.EMIOSPI1SSIN (emio_spi1_ss_i_n),
.EMIOSPI1SSON ({emio_spi1_ss2_o_n,emio_spi1_ss1_o_n,emio_spi1_ss_o_n}),
.EMIOSPI1SSNTN (emio_spi1_ss_n_t_n),
.PLPSTRACECLK (clk_pl_to_ps_trace),
.PSPLTRACECTL (ps_pl_tracectl),
.PSPLTRACEDATA (ps_pl_tracedata),
.EMIOTTC0WAVEO (emio_ttc0_wave_o),
.EMIOTTC0CLKI (clk_pl_to_ps_emio_ttc0),
.EMIOTTC1WAVEO (emio_ttc1_wave_o),
.EMIOTTC1CLKI (clk_pl_to_ps_emio_ttc1),
.EMIOTTC2WAVEO (emio_ttc2_wave_o),
.EMIOTTC2CLKI (clk_pl_to_ps_emio_ttc2),
.EMIOTTC3WAVEO (emio_ttc3_wave_o),
.EMIOTTC3CLKI (clk_pl_to_ps_emio_ttc3),
.EMIOWDT0CLKI (clk_pl_to_ps_emio_wdt0),
.EMIOWDT0RSTO (emio_wdt0_rst_o),
.EMIOWDT1CLKI (clk_pl_to_ps_emio_wdt1),
.EMIOWDT1RSTO (emio_wdt1_rst_o),
.EMIOHUBPORTOVERCRNTUSB30 (emio_hub_port_overcrnt_usb3_0),
.EMIOHUBPORTOVERCRNTUSB31 (emio_hub_port_overcrnt_usb3_1),
.EMIOHUBPORTOVERCRNTUSB20 (emio_hub_port_overcrnt_usb2_0),
.EMIOHUBPORTOVERCRNTUSB21 (emio_hub_port_overcrnt_usb2_1),
.EMIOU2DSPORTVBUSCTRLUSB30 (emio_u2dsport_vbus_ctrl_usb3_0),
.EMIOU2DSPORTVBUSCTRLUSB31 (emio_u2dsport_vbus_ctrl_usb3_1),
.EMIOU3DSPORTVBUSCTRLUSB30 (emio_u3dsport_vbus_ctrl_usb3_0),
.EMIOU3DSPORTVBUSCTRLUSB31 (emio_u3dsport_vbus_ctrl_usb3_1),
.ADMAFCICLK (clk_pl_to_ps_adma_fci),
.PL2ADMACVLD (pl2adma_cvld),
.PL2ADMATACK (pl2adma_tack),
.ADMA2PLCACK (adma2pl_cack),
.ADMA2PLTVLD (adma2pl_tvld),
.GDMAFCICLK (clk_pl_to_ps_gdma_perif),
.PL2GDMACVLD (perif_gdma_cvld),
.PL2GDMATACK (perif_gdma_tack),
.GDMA2PLCACK (gdma_perif_cack),
.GDMA2PLTVLD (gdma_perif_tvld),
.PLFPGASTOP (pl_clock_stop),
.PLLAUXREFCLKLPD (clk_pl_to_ps_pll_aux_lpd),
.PLLAUXREFCLKFPD (clk_pl_to_ps_pll_aux_fpd),
.DPSAXISAUDIOTDATA (pl_to_ps_axi_stream_dp_audio_tdata),
.DPSAXISAUDIOTID (pl_to_ps_axi_stream_dp_audio_tid),
.DPSAXISAUDIOTVALID (pl_to_ps_axi_stream_dp_audio_tvalid),
.DPSAXISAUDIOTREADY (pl_to_ps_axi_stream_dp_audio_tready),
.DPMAXISMIXEDAUDIOTDATA (ps_to_pl_axi_stream_dp_mixed_audio_tdata),
.DPMAXISMIXEDAUDIOTID (ps_to_pl_axi_stream_dp_mixed_audio_tid),
.DPMAXISMIXEDAUDIOTVALID (ps_to_pl_axi_stream_dp_mixed_audio_tvalid),
.DPMAXISMIXEDAUDIOTREADY (ps_to_pl_axi_stream_dp_mixed_audio_tready),
.DPSAXISAUDIOCLK (clk_pl_to_ps_dp_s_axis_audio),
.DPLIVEVIDEOINVSYNC (dp_live_video_in_vsync),
.DPLIVEVIDEOINHSYNC (dp_live_video_in_hsync),
.DPLIVEVIDEOINDE (dp_live_video_in_de),
.DPLIVEVIDEOINPIXEL1 (dp_live_video_in_pixel1),
.DPVIDEOINCLK (clk_pl_to_ps_dp_video_in),
.DPVIDEOOUTHSYNC (dp_video_out_hsync),
.DPVIDEOOUTVSYNC (dp_video_out_vsync),
.DPVIDEOOUTPIXEL1 (dp_video_out_pixel1),
.DPAUXDATAIN (dp_aux_data_in),
.DPAUXDATAOUT (dp_aux_data_out),
.DPAUXDATAOEN (dp_aux_data_oe_n),
.DPLIVEGFXALPHAIN (dp_live_gfx_alpha_in),
.DPLIVEGFXPIXEL1IN (dp_live_gfx_pixel1_in),
.DPHOTPLUGDETECT (dp_hot_plug_detect),
.DPEXTERNALCUSTOMEVENT1 (dp_external_custom_event1),
.DPEXTERNALCUSTOMEVENT2 (dp_external_custom_event2),
.DPEXTERNALVSYNCEVENT (dp_external_vsync_event),
.DPLIVEVIDEODEOUT (dp_live_video_de_out),
.PLPSEVENTI (pl_ps_eventi),
.PSPLEVENTO (ps_pl_evento),
.PSPLSTANDBYWFE (ps_pl_standbywfe),
.PSPLSTANDBYWFI (ps_pl_standbywfi),
.PLPSAPUGICIRQ (pl_ps_apugic_irq),
.PLPSAPUGICFIQ (pl_ps_apugic_fiq),
.RPUEVENTI0 (rpu_eventi0),
.RPUEVENTI1 (rpu_eventi1),
.RPUEVENTO0 (rpu_evento0),
.RPUEVENTO1 (rpu_evento1),
.NFIQ0LPDRPU (nfiq0_lpd_rpu),
.NFIQ1LPDRPU (nfiq1_lpd_rpu),
.NIRQ0LPDRPU (nirq0_lpd_rpu),
.NIRQ1LPDRPU (nirq1_lpd_rpu),
.STMEVENT (stm_event),
.PLPSTRIGACK (pl_ps_trigack),
.PLPSTRIGGER (pl_ps_trigger),
.PSPLTRIGACK (ps_pl_trigack),
.PSPLTRIGGER (ps_pl_trigger),
.FTMGPO (ftm_gpo),
.FTMGPI (ftm_gpi),
.PLPSIRQ0 (pl_ps_irq0),
.PLPSIRQ1 (pl_ps_irq1),
.PSPLIRQLPD ({irq_lpd_dev_null[18:8],
							ps_to_pl_irq_xmpu_lpd,
							ps_to_pl_irq_efuse,
							ps_to_pl_irq_csu_dma,
							ps_to_pl_irq_csu,
							ps_to_pl_irq_adma_chan,
							ps_to_pl_irq_usb3_0_pmu_wakeup,
							ps_to_pl_irq_usb3_1_otg,
							ps_to_pl_irq_usb3_1_endpoint,
							ps_to_pl_irq_usb3_0_otg,
							ps_to_pl_irq_usb3_0_endpoint,
							ps_to_pl_irq_enet3_wake,
							ps_to_pl_irq_enet3,
							ps_to_pl_irq_enet2_wake,
							ps_to_pl_irq_enet2,
							ps_to_pl_irq_enet1_wake,
							ps_to_pl_irq_enet1,
							ps_to_pl_irq_enet0_wake,
							ps_to_pl_irq_enet0,
							ps_to_pl_irq_ams,
							ps_to_pl_irq_aib_axi,
							ps_to_pl_irq_atb_err_lpd,
							ps_to_pl_irq_csu_pmu_wdt,
							ps_to_pl_irq_lp_wdt,
							ps_to_pl_irq_sdio1_wake,
							ps_to_pl_irq_sdio0_wake,
							ps_to_pl_irq_sdio1,
							ps_to_pl_irq_sdio0,
							ps_to_pl_irq_ttc3_2,
							ps_to_pl_irq_ttc3_1,
							ps_to_pl_irq_ttc3_0,
							ps_to_pl_irq_ttc2_2,
							ps_to_pl_irq_ttc2_1,
							ps_to_pl_irq_ttc2_0,
							ps_to_pl_irq_ttc1_2,
							ps_to_pl_irq_ttc1_1,
							ps_to_pl_irq_ttc1_0,
							ps_to_pl_irq_ttc0_2,
							ps_to_pl_irq_ttc0_1,
							ps_to_pl_irq_ttc0_0,
							ps_to_pl_irq_ipi_channel0,
							ps_to_pl_irq_ipi_channel1,
							ps_to_pl_irq_ipi_channel2,
							ps_to_pl_irq_ipi_channel7,
							ps_to_pl_irq_ipi_channel8,
							ps_to_pl_irq_ipi_channel9,
							ps_to_pl_irq_ipi_channel10,
							ps_to_pl_irq_clkmon,
							ps_to_pl_irq_rtc_seconds,
							ps_to_pl_irq_rtc_alaram,
							ps_to_pl_irq_lpd_apm,
							ps_to_pl_irq_can1,
							ps_to_pl_irq_can0,
							ps_to_pl_irq_uart1,
							ps_to_pl_irq_uart0,
							ps_to_pl_irq_spi1,
							ps_to_pl_irq_spi0,
							ps_to_pl_irq_i2c1,
							ps_to_pl_irq_i2c0,
							ps_to_pl_irq_gpio,
							ps_to_pl_irq_qspi,
							ps_to_pl_irq_nand,
							ps_to_pl_irq_r5_core1_ecc_error,
							ps_to_pl_irq_r5_core0_ecc_error,
							ps_to_pl_irq_lpd_apb_intr,
							ps_to_pl_irq_ocm_error,
							ps_to_pl_irq_rpu_pm,
							irq_lpd_dev_null[7:0]}),
.PSPLIRQFPD ({irq_fpd_dev_null[19:12],
							ps_to_pl_irq_intf_fpd_smmu,
							ps_to_pl_irq_intf_ppd_cci,
							ps_to_pl_irq_apu_regs,
							ps_to_pl_irq_apu_exterr,
							ps_to_pl_irq_apu_l2err,
							ps_to_pl_irq_apu_comm,
							ps_to_pl_irq_apu_pmu,
							ps_to_pl_irq_apu_cti,
							ps_to_pl_irq_apu_cpumnt,
							ps_to_pl_irq_xmpu_fpd,
							ps_to_pl_irq_sata,
							ps_to_pl_irq_gpu,
							ps_to_pl_irq_gdma_chan,
							ps_to_pl_irq_apm_fpd,
							ps_to_pl_irq_dpdma,
							ps_to_pl_irq_fpd_atb_error,
							ps_to_pl_irq_fpd_apb_int,
							ps_to_pl_irq_dport,
							ps_to_pl_irq_pcie_msc,
							ps_to_pl_irq_pcie_dma,
							ps_to_pl_irq_pcie_legacy,
							ps_to_pl_irq_pcie_msi,
							ps_to_pl_irq_fp_wdt,
							ps_to_pl_irq_ddr_ss,
							irq_fpd_dev_null[11:0]}),
.OSCRTCCLK (osc_rtc_clk),
.PLPMUGPI (pl_pmu_gpi),
.PMUPLGPO (pmu_pl_gpo),
.AIBPMUAFIFMFPDACK (aib_pmu_afifm_fpd_ack),
.AIBPMUAFIFMLPDACK (aib_pmu_afifm_lpd_ack),
.PMUAIBAFIFMFPDREQ (pmu_aib_afifm_fpd_req),
.PMUAIBAFIFMLPDREQ (pmu_aib_afifm_lpd_req),
.PMUERRORTOPL (pmu_error_to_pl),
.PMUERRORFROMPL (pmu_error_from_pl),
.DDRCEXTREFRESHRANK0REQ (ddrc_ext_refresh_rank0_req),
.DDRCEXTREFRESHRANK1REQ (ddrc_ext_refresh_rank1_req),
.DDRCREFRESHPLCLK (clk_pl_to_ps_ddrc_refresh),
.PLACPINACT (pl_acpinact),
.PLCLK (clk_ps_to_pl_clks),
.DPVIDEOREFCLK(clk_ps_to_pl_dp_video),
.DPAUDIOREFCLK(clk_ps_to_pl_dp_audio),
.PSS_ALTO_CORE_PAD_MGTTXN0OUT(pss_alto_core_pad_mgttxn0out),// What are these?
.PSS_ALTO_CORE_PAD_MGTTXN1OUT(pss_alto_core_pad_mgttxn1out),
.PSS_ALTO_CORE_PAD_MGTTXN2OUT(pss_alto_core_pad_mgttxn2out),
.PSS_ALTO_CORE_PAD_MGTTXN3OUT(pss_alto_core_pad_mgttxn3out),
.PSS_ALTO_CORE_PAD_MGTTXP0OUT(pss_alto_core_pad_mgttxp0out),
.PSS_ALTO_CORE_PAD_MGTTXP1OUT(pss_alto_core_pad_mgttxp1out),
.PSS_ALTO_CORE_PAD_MGTTXP2OUT(pss_alto_core_pad_mgttxp2out),
.PSS_ALTO_CORE_PAD_MGTTXP3OUT(pss_alto_core_pad_mgttxp3out),
.PSS_ALTO_CORE_PAD_PADO(pss_alto_core_pad_pad0),
.PSS_ALTO_CORE_PAD_BOOTMODE(),
.PSS_ALTO_CORE_PAD_CLK(),
.PSS_ALTO_CORE_PAD_DONEB(),
.PSS_ALTO_CORE_PAD_DRAMA(),
.PSS_ALTO_CORE_PAD_DRAMACTN(),
.PSS_ALTO_CORE_PAD_DRAMALERTN(),
.PSS_ALTO_CORE_PAD_DRAMBA(),
.PSS_ALTO_CORE_PAD_DRAMBG(),
.PSS_ALTO_CORE_PAD_DRAMCK(),
.PSS_ALTO_CORE_PAD_DRAMCKE(),
.PSS_ALTO_CORE_PAD_DRAMCKN(),
.PSS_ALTO_CORE_PAD_DRAMCSN(),
.PSS_ALTO_CORE_PAD_DRAMDM(),
.PSS_ALTO_CORE_PAD_DRAMDQ(),
.PSS_ALTO_CORE_PAD_DRAMDQS(),
.PSS_ALTO_CORE_PAD_DRAMDQSN(),
.PSS_ALTO_CORE_PAD_DRAMODT(),
.PSS_ALTO_CORE_PAD_DRAMPARITY(),
.PSS_ALTO_CORE_PAD_DRAMRAMRSTN(),
.PSS_ALTO_CORE_PAD_ERROROUT(),
.PSS_ALTO_CORE_PAD_ERRORSTATUS(),
.PSS_ALTO_CORE_PAD_INITB(),
.PSS_ALTO_CORE_PAD_JTAGTCK(),
.PSS_ALTO_CORE_PAD_JTAGTDI(),
.PSS_ALTO_CORE_PAD_JTAGTDO(),
.PSS_ALTO_CORE_PAD_JTAGTMS(),
.PSS_ALTO_CORE_PAD_MIO(),
.PSS_ALTO_CORE_PAD_PORB(),
.PSS_ALTO_CORE_PAD_PROGB(),
.PSS_ALTO_CORE_PAD_RCALIBINOUT(),
.PSS_ALTO_CORE_PAD_SRSTB(),
.PSS_ALTO_CORE_PAD_ZQ(),
.PSS_ALTO_CORE_PAD_MGTRXN0IN(),
.PSS_ALTO_CORE_PAD_MGTRXN1IN(),
.PSS_ALTO_CORE_PAD_MGTRXN2IN(),
.PSS_ALTO_CORE_PAD_MGTRXN3IN(),
.PSS_ALTO_CORE_PAD_MGTRXP0IN(),
.PSS_ALTO_CORE_PAD_MGTRXP1IN(),
.PSS_ALTO_CORE_PAD_MGTRXP2IN(),
.PSS_ALTO_CORE_PAD_MGTRXP3IN(),
.PSS_ALTO_CORE_PAD_PADI(),
.PSS_ALTO_CORE_PAD_REFN0IN(),
.PSS_ALTO_CORE_PAD_REFN1IN(),
.PSS_ALTO_CORE_PAD_REFN2IN(),
.PSS_ALTO_CORE_PAD_REFN3IN(),
.PSS_ALTO_CORE_PAD_REFP0IN(),
.PSS_ALTO_CORE_PAD_REFP1IN(),
.PSS_ALTO_CORE_PAD_REFP2IN(),
.PSS_ALTO_CORE_PAD_REFP3IN()
);

endmodule
