// [5:0]AxUSER driven by PL-AXI_ID
// [15:6]AxUSER need to be tied to 10'b0000001111

module RawPS8(

// Clocks (all unbuffered)
// from ps to pl (fps_tpl)
output wire clk_fps_tpl_dp_video,
output wire clk_fps_tpl_dp_audio,
output wire clk_fps_tpl_fmio_gem0_fifo_tx,
output wire clk_fps_tpl_fmio_gem0_fifo_rx,
output wire clk_fps_tpl_fmio_gem1_fifo_tx,
output wire clk_fps_tpl_fmio_gem1_fifo_rx,
output wire clk_fps_tpl_fmio_gem2_fifo_tx,
output wire clk_fps_tpl_fmio_gem2_fifo_rx,
output wire clk_fps_tpl_fmio_gem3_fifo_tx,
output wire clk_fps_tpl_fmio_gem3_fifo_rx,
output wire clk_fps_tpl_gem_tsu_clk,
output wire clk_fps_tpl_emio_sdio0,
output wire clk_fps_tpl_emio_sdio1,
output wire clk_fps_tpl_trace,
output wire [3:0] clk_fps_tpl_clks,

// to ps from pl (tps_fpl)
input  wire clk_tps_fpl_supplier_axi_hpm0_fpd, // dp + supplier gp0
input  wire clk_tps_fpl_supplier_axi_hpm0_lpd, // supplier gp2
input  wire clk_tps_fpl_supplier_axi_hpm1_fpd, // supplier gp1
input  wire clk_tps_fpl_consumer_axi_hpc0_fpd_read,  // consumer gp0 read
input  wire clk_tps_fpl_consumer_axi_hpc0_fpd_write, // consumer gp0 write
input  wire clk_tps_fpl_consumer_axi_hpc1_fpd_read,  // consumer gp1 read
input  wire clk_tps_fpl_consumer_axi_hpc1_fpd_write, // consumer gp1 write
input  wire clk_tps_fpl_consumer_axi_hp0_fpd_read,   // consumer gp2 read
input  wire clk_tps_fpl_consumer_axi_hp0_fpd_write,  // consumer gp2 write
input  wire clk_tps_fpl_consumer_axi_hp1_fpd_read,   // consumer gp3 read
input  wire clk_tps_fpl_consumer_axi_hp1_fpd_write,  // consumer gp3 write
input  wire clk_tps_fpl_consumer_axi_hp2_fpd_read,   // consumer gp4 read
input  wire clk_tps_fpl_consumer_axi_hp2_fpd_write,  // consumer gp4 write
input  wire clk_tps_fpl_consumer_axi_hp3_fpd_read,   // consumer gp5 read
input  wire clk_tps_fpl_consumer_axi_hp3_fpd_write,  // consumer gp5 write
input  wire clk_tps_fpl_consumer_axi_lpd_read,       // consumer gp6 read
input  wire clk_tps_fpl_consumer_axi_lpd_write,      // consumer gp6 write
input  wire clk_tps_fpl_consumer_axi_acp_fpd,            // consumer acp
input  wire clk_tps_fpl_consumer_axi_ace_fpd,            // consumer ace
input  wire clk_tps_fpl_emio_enet0_gmii_rx,
input  wire clk_tps_fpl_emio_enet0_gmii_tx,
input  wire clk_tps_fpl_emio_enet1_gmii_rx,
input  wire clk_tps_fpl_emio_enet1_gmii_tx,
input  wire clk_tps_fpl_emio_enet2_gmii_rx,
input  wire clk_tps_fpl_emio_enet2_gmii_tx,
input  wire clk_tps_fpl_emio_enet3_gmii_rx,
input  wire clk_tps_fpl_emio_enet3_gmii_tx,
input wire  clk_tps_fpl_fmio_gem0_fifo_tx,
input wire  clk_tps_fpl_fmio_gem0_fifo_rx,
input wire  clk_tps_fpl_fmio_gem1_fifo_tx,
input wire  clk_tps_fpl_fmio_gem1_fifo_rx,
input wire  clk_tps_fpl_fmio_gem2_fifo_tx,
input wire  clk_tps_fpl_fmio_gem2_fifo_rx,
input wire  clk_tps_fpl_fmio_gem3_fifo_tx,
input wire  clk_tps_fpl_fmio_gem3_fifo_rx,
input wire  clk_tps_fpl_fmio_gem_tsu,
input  wire clk_tps_fpl_emio_enet_tsu,
input  wire clk_tps_fpl_emio_sdio0,
input  wire clk_tps_fpl_emio_sdio1,     
input wire clk_tps_fpl_trace,
input  wire [2:0] clk_tps_fpl_emio_ttc0,
input  wire [2:0] clk_tps_fpl_emio_ttc1,
input  wire [2:0] clk_tps_fpl_emio_ttc2,
input  wire [2:0] clk_tps_fpl_emio_ttc3,
input  wire clk_tps_fpl_emio_wdt0,
input  wire clk_tps_fpl_emio_wdt1,
input  wire [7:0] clk_tps_fpl_adma_fci,
input  wire [7:0] clk_tps_fpl_gdma_perif,
input  wire [1:0] clk_tps_fpl_pll_aux_lpd,
input  wire [2:0] clk_tps_fpl_pll_aux_fpd,
input  wire clk_tps_fpl_dp_s_axis_audio,
input  wire clk_tps_fpl_dp_video_in,
input  wire clk_tps_fpl_ddrc_refresh,
input  [3:0]  clk_tps_fpl_pstp,

// axi interfaces ports
// 3 128 bit supplier axi interfaces
// 8 128 bit consumer axi interfaces
output wire [15:0]   supplier_axi_gp0_awid,
output wire [39:0]   supplier_axi_gp0_awaddr, 
output wire [7:0]    supplier_axi_gp0_awlen,  
output wire [2:0]    supplier_axi_gp0_awsize, 
output wire [1:0]    supplier_axi_gp0_awburst,
output wire          supplier_axi_gp0_awlock, 
output wire [3:0]    supplier_axi_gp0_awcache,
output wire [2:0]    supplier_axi_gp0_awprot, 
output wire          supplier_axi_gp0_awvalid,
output wire [15:0]   supplier_axi_gp0_awuser, 
input  wire          supplier_axi_gp0_awready,
output wire [127:0]  supplier_axi_gp0_wdata,  
output wire [15:0]   supplier_axi_gp0_wstrb,  
output wire          supplier_axi_gp0_wlast,  
output wire          supplier_axi_gp0_wvalid, 
input  wire          supplier_axi_gp0_wready, 
input  wire [15:0]   supplier_axi_gp0_bid,    
input  wire [1:0]    supplier_axi_gp0_bresp,  
input  wire          supplier_axi_gp0_bvalid, 
output wire          supplier_axi_gp0_bready, 
output wire [15:0]   supplier_axi_gp0_arid,   
output wire [39:0]   supplier_axi_gp0_araddr, 
output wire [7:0]    supplier_axi_gp0_arlen,  
output wire [2:0]    supplier_axi_gp0_arsize, 
output wire [1:0]    supplier_axi_gp0_arburst,
output wire          supplier_axi_gp0_arlock, 
output wire [3:0]    supplier_axi_gp0_arcache,
output wire [2:0]    supplier_axi_gp0_arprot, 
output wire          supplier_axi_gp0_arvalid,
output wire [15:0]   supplier_axi_gp0_aruser, 
input  wire          supplier_axi_gp0_arready,
input  wire [15:0]   supplier_axi_gp0_rid,    
input  wire [127:0]  supplier_axi_gp0_rdata,  
input  wire [1:0]    supplier_axi_gp0_rresp,  
input  wire          supplier_axi_gp0_rlast,  
input  wire          supplier_axi_gp0_rvalid, 
output wire          supplier_axi_gp0_rready, 
output wire [3:0]    supplier_axi_gp0_awqos,  
output wire [3:0]    supplier_axi_gp0_arqos,  

output wire [15:0]   supplier_axi_gp1_awid,
output wire [39:0]   supplier_axi_gp1_awaddr, 
output wire [7:0]    supplier_axi_gp1_awlen,  
output wire [2:0]    supplier_axi_gp1_awsize, 
output wire [1:0]    supplier_axi_gp1_awburst,
output wire          supplier_axi_gp1_awlock, 
output wire [3:0]    supplier_axi_gp1_awcache,
output wire [2:0]    supplier_axi_gp1_awprot, 
output wire          supplier_axi_gp1_awvalid,
output wire [15:0]   supplier_axi_gp1_awuser, 
input  wire          supplier_axi_gp1_awready,
output wire [127:0]  supplier_axi_gp1_wdata,  
output wire [15:0]   supplier_axi_gp1_wstrb,  
output wire          supplier_axi_gp1_wlast,  
output wire          supplier_axi_gp1_wvalid, 
input  wire          supplier_axi_gp1_wready, 
input  wire [15:0]   supplier_axi_gp1_bid,    
input  wire [1:0]    supplier_axi_gp1_bresp,  
input  wire          supplier_axi_gp1_bvalid, 
output wire          supplier_axi_gp1_bready, 
output wire [15:0]   supplier_axi_gp1_arid,   
output wire [39:0]   supplier_axi_gp1_araddr, 
output wire [7:0]    supplier_axi_gp1_arlen,  
output wire [2:0]    supplier_axi_gp1_arsize, 
output wire [1:0]    supplier_axi_gp1_arburst,
output wire          supplier_axi_gp1_arlock, 
output wire [3:0]    supplier_axi_gp1_arcache,
output wire [2:0]    supplier_axi_gp1_arprot, 
output wire          supplier_axi_gp1_arvalid,
output wire [15:0]   supplier_axi_gp1_aruser, 
input  wire          supplier_axi_gp1_arready,
input  wire [15:0]   supplier_axi_gp1_rid,    
input  wire [127:0]  supplier_axi_gp1_rdata,  
input  wire [1:0]    supplier_axi_gp1_rresp,  
input  wire          supplier_axi_gp1_rlast,  
input  wire          supplier_axi_gp1_rvalid, 
output wire          supplier_axi_gp1_rready, 
output wire [3:0]    supplier_axi_gp1_awqos,  
output wire [3:0]    supplier_axi_gp1_arqos,  

output wire [15:0]   supplier_axi_gp2_awid,
output wire [39:0]   supplier_axi_gp2_awaddr, 
output wire [7:0]    supplier_axi_gp2_awlen,  
output wire [2:0]    supplier_axi_gp2_awsize, 
output wire [1:0]    supplier_axi_gp2_awburst,
output wire          supplier_axi_gp2_awlock, 
output wire [3:0]    supplier_axi_gp2_awcache,
output wire [2:0]    supplier_axi_gp2_awprot, 
output wire          supplier_axi_gp2_awvalid,
output wire [15:0]   supplier_axi_gp2_awuser, 
input  wire          supplier_axi_gp2_awready,
output wire [127:0]  supplier_axi_gp2_wdata,  
output wire [15:0]   supplier_axi_gp2_wstrb,  
output wire          supplier_axi_gp2_wlast,  
output wire          supplier_axi_gp2_wvalid, 
input  wire          supplier_axi_gp2_wready, 
input  wire [15:0]   supplier_axi_gp2_bid,    
input  wire [1:0]    supplier_axi_gp2_bresp,  
input  wire          supplier_axi_gp2_bvalid, 
output wire          supplier_axi_gp2_bready, 
output wire [15:0]   supplier_axi_gp2_arid,   
output wire [39:0]   supplier_axi_gp2_araddr, 
output wire [7:0]    supplier_axi_gp2_arlen,  
output wire [2:0]    supplier_axi_gp2_arsize, 
output wire [1:0]    supplier_axi_gp2_arburst,
output wire          supplier_axi_gp2_arlock, 
output wire [3:0]    supplier_axi_gp2_arcache,
output wire [2:0]    supplier_axi_gp2_arprot, 
output wire          supplier_axi_gp2_arvalid,
output wire [15:0]   supplier_axi_gp2_aruser, 
input  wire          supplier_axi_gp2_arready,
input  wire [15:0]   supplier_axi_gp2_rid,    
input  wire [127:0]  supplier_axi_gp2_rdata,  
input  wire [1:0]    supplier_axi_gp2_rresp,  
input  wire          supplier_axi_gp2_rlast,  
input  wire          supplier_axi_gp2_rvalid, 
output wire          supplier_axi_gp2_rready, 
output wire [3:0]    supplier_axi_gp2_awqos,  
output wire [3:0]    supplier_axi_gp2_arqos,  

input  wire          consumer_axi_gp0_aruser,
input  wire          consumer_axi_gp0_awuser, 
input  wire [5:0]    consumer_axi_gp0_awid,   
input  wire [48:0]   consumer_axi_gp0_awaddr, 
input  wire [7:0]    consumer_axi_gp0_awlen , 
input  wire [2:0]    consumer_axi_gp0_awsize, 
input  wire [1:0]    consumer_axi_gp0_awburst,
input  wire          consumer_axi_gp0_awlock, 
input  wire [3:0]    consumer_axi_gp0_awcache,
input  wire [2:0]    consumer_axi_gp0_awprot, 
input  wire          consumer_axi_gp0_awvalid,
output wire          consumer_axi_gp0_awready,
input  wire [127:0]  consumer_axi_gp0_wdata,  
input  wire [15:0]   consumer_axi_gp0_wstrb, 
input  wire          consumer_axi_gp0_wlast,  
input  wire          consumer_axi_gp0_wvalid, 
output wire          consumer_axi_gp0_wready, 
output wire [5:0]    consumer_axi_gp0_bid,    
output wire [1:0]    consumer_axi_gp0_bresp,  
output wire          consumer_axi_gp0_bvalid, 
input  wire          consumer_axi_gp0_bready, 
input  wire [5:0]    consumer_axi_gp0_arid,   
input  wire [48:0]   consumer_axi_gp0_araddr, 
input  wire [7:0]    consumer_axi_gp0_arlen,  
input  wire [2:0]    consumer_axi_gp0_arsize, 
input  wire [1:0]    consumer_axi_gp0_arburst,
input  wire          consumer_axi_gp0_arlock, 
input  wire [3:0]    consumer_axi_gp0_arcache,
input  wire [2:0]    consumer_axi_gp0_arprot, 
input  wire          consumer_axi_gp0_arvalid,
output wire          consumer_axi_gp0_arready,
output wire [5:0]    consumer_axi_gp0_rid,    
output wire [127:0]  consumer_axi_gp0_rdata,  
output wire [1:0]    consumer_axi_gp0_rresp,  
output wire          consumer_axi_gp0_rlast,  
output wire          consumer_axi_gp0_rvalid, 
input  wire          consumer_axi_gp0_rready, 
input  wire [3:0]    consumer_axi_gp0_awqos,  
input  wire [3:0]    consumer_axi_gp0_arqos,  
output wire [7:0]    consumer_axi_gp0_rcount, 
output wire [7:0]    consumer_axi_gp0_wcount, 
output wire [3:0]    consumer_axi_gp0_racount,
output wire [3:0]    consumer_axi_gp0_wacount,

input  wire          consumer_axi_gp1_aruser,
input  wire          consumer_axi_gp1_awuser, 
input  wire [5:0]    consumer_axi_gp1_awid,   
input  wire [48:0]   consumer_axi_gp1_awaddr, 
input  wire [7:0]    consumer_axi_gp1_awlen , 
input  wire [2:0]    consumer_axi_gp1_awsize, 
input  wire [1:0]    consumer_axi_gp1_awburst,
input  wire          consumer_axi_gp1_awlock, 
input  wire [3:0]    consumer_axi_gp1_awcache,
input  wire [2:0]    consumer_axi_gp1_awprot, 
input  wire          consumer_axi_gp1_awvalid,
output wire          consumer_axi_gp1_awready,
input  wire [127:0]  consumer_axi_gp1_wdata,  
input  wire [15:0]   consumer_axi_gp1_wstrb, 
input  wire          consumer_axi_gp1_wlast,  
input  wire          consumer_axi_gp1_wvalid, 
output wire          consumer_axi_gp1_wready, 
output wire [5:0]    consumer_axi_gp1_bid,    
output wire [1:0]    consumer_axi_gp1_bresp,  
output wire          consumer_axi_gp1_bvalid, 
input  wire          consumer_axi_gp1_bready, 
input  wire [5:0]    consumer_axi_gp1_arid,   
input  wire [48:0]   consumer_axi_gp1_araddr, 
input  wire [7:0]    consumer_axi_gp1_arlen,  
input  wire [2:0]    consumer_axi_gp1_arsize, 
input  wire [1:0]    consumer_axi_gp1_arburst,
input  wire          consumer_axi_gp1_arlock, 
input  wire [3:0]    consumer_axi_gp1_arcache,
input  wire [2:0]    consumer_axi_gp1_arprot, 
input  wire          consumer_axi_gp1_arvalid,
output wire          consumer_axi_gp1_arready,
output wire [5:0]    consumer_axi_gp1_rid,    
output wire [127:0]  consumer_axi_gp1_rdata,  
output wire [1:0]    consumer_axi_gp1_rresp,  
output wire          consumer_axi_gp1_rlast,  
output wire          consumer_axi_gp1_rvalid, 
input  wire          consumer_axi_gp1_rready, 
input  wire [3:0]    consumer_axi_gp1_awqos,  
input  wire [3:0]    consumer_axi_gp1_arqos,  
output wire [7:0]    consumer_axi_gp1_rcount, 
output wire [7:0]    consumer_axi_gp1_wcount, 
output wire [3:0]    consumer_axi_gp1_racount,
output wire [3:0]    consumer_axi_gp1_wacount,

input  wire          consumer_axi_gp2_aruser,
input  wire          consumer_axi_gp2_awuser, 
input  wire [5:0]    consumer_axi_gp2_awid,   
input  wire [48:0]   consumer_axi_gp2_awaddr, 
input  wire [7:0]    consumer_axi_gp2_awlen , 
input  wire [2:0]    consumer_axi_gp2_awsize, 
input  wire [1:0]    consumer_axi_gp2_awburst,
input  wire          consumer_axi_gp2_awlock, 
input  wire [3:0]    consumer_axi_gp2_awcache,
input  wire [2:0]    consumer_axi_gp2_awprot, 
input  wire          consumer_axi_gp2_awvalid,
output wire          consumer_axi_gp2_awready,
input  wire [127:0]  consumer_axi_gp2_wdata,  
input  wire [15:0]   consumer_axi_gp2_wstrb, 
input  wire          consumer_axi_gp2_wlast,  
input  wire          consumer_axi_gp2_wvalid, 
output wire          consumer_axi_gp2_wready, 
output wire [5:0]    consumer_axi_gp2_bid,    
output wire [1:0]    consumer_axi_gp2_bresp,  
output wire          consumer_axi_gp2_bvalid, 
input  wire          consumer_axi_gp2_bready, 
input  wire [5:0]    consumer_axi_gp2_arid,   
input  wire [48:0]   consumer_axi_gp2_araddr, 
input  wire [7:0]    consumer_axi_gp2_arlen,  
input  wire [2:0]    consumer_axi_gp2_arsize, 
input  wire [1:0]    consumer_axi_gp2_arburst,
input  wire          consumer_axi_gp2_arlock, 
input  wire [3:0]    consumer_axi_gp2_arcache,
input  wire [2:0]    consumer_axi_gp2_arprot, 
input  wire          consumer_axi_gp2_arvalid,
output wire          consumer_axi_gp2_arready,
output wire [5:0]    consumer_axi_gp2_rid,    
output wire [127:0]  consumer_axi_gp2_rdata,  
output wire [1:0]    consumer_axi_gp2_rresp,  
output wire          consumer_axi_gp2_rlast,  
output wire          consumer_axi_gp2_rvalid, 
input  wire          consumer_axi_gp2_rready, 
input  wire [3:0]    consumer_axi_gp2_awqos,  
input  wire [3:0]    consumer_axi_gp2_arqos,  
output wire [7:0]    consumer_axi_gp2_rcount, 
output wire [7:0]    consumer_axi_gp2_wcount, 
output wire [3:0]    consumer_axi_gp2_racount,
output wire [3:0]    consumer_axi_gp2_wacount,

input  wire          consumer_axi_gp3_aruser,
input  wire          consumer_axi_gp3_awuser, 
input  wire [5:0]    consumer_axi_gp3_awid,   
input  wire [48:0]   consumer_axi_gp3_awaddr, 
input  wire [7:0]    consumer_axi_gp3_awlen , 
input  wire [2:0]    consumer_axi_gp3_awsize, 
input  wire [1:0]    consumer_axi_gp3_awburst,
input  wire          consumer_axi_gp3_awlock, 
input  wire [3:0]    consumer_axi_gp3_awcache,
input  wire [2:0]    consumer_axi_gp3_awprot, 
input  wire          consumer_axi_gp3_awvalid,
output wire          consumer_axi_gp3_awready,
input  wire [127:0]  consumer_axi_gp3_wdata,  
input  wire [15:0]   consumer_axi_gp3_wstrb, 
input  wire          consumer_axi_gp3_wlast,  
input  wire          consumer_axi_gp3_wvalid, 
output wire          consumer_axi_gp3_wready, 
output wire [5:0]    consumer_axi_gp3_bid,    
output wire [1:0]    consumer_axi_gp3_bresp,  
output wire          consumer_axi_gp3_bvalid, 
input  wire          consumer_axi_gp3_bready, 
input  wire [5:0]    consumer_axi_gp3_arid,   
input  wire [48:0]   consumer_axi_gp3_araddr, 
input  wire [7:0]    consumer_axi_gp3_arlen,  
input  wire [2:0]    consumer_axi_gp3_arsize, 
input  wire [1:0]    consumer_axi_gp3_arburst,
input  wire          consumer_axi_gp3_arlock, 
input  wire [3:0]    consumer_axi_gp3_arcache,
input  wire [2:0]    consumer_axi_gp3_arprot, 
input  wire          consumer_axi_gp3_arvalid,
output wire          consumer_axi_gp3_arready,
output wire [5:0]    consumer_axi_gp3_rid,    
output wire [127:0]  consumer_axi_gp3_rdata,  
output wire [1:0]    consumer_axi_gp3_rresp,  
output wire          consumer_axi_gp3_rlast,  
output wire          consumer_axi_gp3_rvalid, 
input  wire          consumer_axi_gp3_rready, 
input  wire [3:0]    consumer_axi_gp3_awqos,  
input  wire [3:0]    consumer_axi_gp3_arqos,  
output wire [7:0]    consumer_axi_gp3_rcount, 
output wire [7:0]    consumer_axi_gp3_wcount, 
output wire [3:0]    consumer_axi_gp3_racount,
output wire [3:0]    consumer_axi_gp3_wacount,

input  wire          consumer_axi_gp4_aruser,
input  wire          consumer_axi_gp4_awuser, 
input  wire [5:0]    consumer_axi_gp4_awid,   
input  wire [48:0]   consumer_axi_gp4_awaddr, 
input  wire [7:0]    consumer_axi_gp4_awlen , 
input  wire [2:0]    consumer_axi_gp4_awsize, 
input  wire [1:0]    consumer_axi_gp4_awburst,
input  wire          consumer_axi_gp4_awlock, 
input  wire [3:0]    consumer_axi_gp4_awcache,
input  wire [2:0]    consumer_axi_gp4_awprot, 
input  wire          consumer_axi_gp4_awvalid,
output wire          consumer_axi_gp4_awready,
input  wire [127:0]  consumer_axi_gp4_wdata,  
input  wire [15:0]   consumer_axi_gp4_wstrb, 
input  wire          consumer_axi_gp4_wlast,  
input  wire          consumer_axi_gp4_wvalid, 
output wire          consumer_axi_gp4_wready, 
output wire [5:0]    consumer_axi_gp4_bid,    
output wire [1:0]    consumer_axi_gp4_bresp,  
output wire          consumer_axi_gp4_bvalid, 
input  wire          consumer_axi_gp4_bready, 
input  wire [5:0]    consumer_axi_gp4_arid,   
input  wire [48:0]   consumer_axi_gp4_araddr, 
input  wire [7:0]    consumer_axi_gp4_arlen,  
input  wire [2:0]    consumer_axi_gp4_arsize, 
input  wire [1:0]    consumer_axi_gp4_arburst,
input  wire          consumer_axi_gp4_arlock, 
input  wire [3:0]    consumer_axi_gp4_arcache,
input  wire [2:0]    consumer_axi_gp4_arprot, 
input  wire          consumer_axi_gp4_arvalid,
output wire          consumer_axi_gp4_arready,
output wire [5:0]    consumer_axi_gp4_rid,    
output wire [127:0]  consumer_axi_gp4_rdata,  
output wire [1:0]    consumer_axi_gp4_rresp,  
output wire          consumer_axi_gp4_rlast,  
output wire          consumer_axi_gp4_rvalid, 
input  wire          consumer_axi_gp4_rready, 
input  wire [3:0]    consumer_axi_gp4_awqos,  
input  wire [3:0]    consumer_axi_gp4_arqos,  
output wire [7:0]    consumer_axi_gp4_rcount, 
output wire [7:0]    consumer_axi_gp4_wcount, 
output wire [3:0]    consumer_axi_gp4_racount,
output wire [3:0]    consumer_axi_gp4_wacount,

input  wire          consumer_axi_gp5_aruser,
input  wire          consumer_axi_gp5_awuser, 
input  wire [5:0]    consumer_axi_gp5_awid,   
input  wire [48:0]   consumer_axi_gp5_awaddr, 
input  wire [7:0]    consumer_axi_gp5_awlen , 
input  wire [2:0]    consumer_axi_gp5_awsize, 
input  wire [1:0]    consumer_axi_gp5_awburst,
input  wire          consumer_axi_gp5_awlock, 
input  wire [3:0]    consumer_axi_gp5_awcache,
input  wire [2:0]    consumer_axi_gp5_awprot, 
input  wire          consumer_axi_gp5_awvalid,
output wire          consumer_axi_gp5_awready,
input  wire [127:0]  consumer_axi_gp5_wdata,  
input  wire [15:0]   consumer_axi_gp5_wstrb, 
input  wire          consumer_axi_gp5_wlast,  
input  wire          consumer_axi_gp5_wvalid, 
output wire          consumer_axi_gp5_wready, 
output wire [5:0]    consumer_axi_gp5_bid,    
output wire [1:0]    consumer_axi_gp5_bresp,  
output wire          consumer_axi_gp5_bvalid, 
input  wire          consumer_axi_gp5_bready, 
input  wire [5:0]    consumer_axi_gp5_arid,   
input  wire [48:0]   consumer_axi_gp5_araddr, 
input  wire [7:0]    consumer_axi_gp5_arlen,  
input  wire [2:0]    consumer_axi_gp5_arsize, 
input  wire [1:0]    consumer_axi_gp5_arburst,
input  wire          consumer_axi_gp5_arlock, 
input  wire [3:0]    consumer_axi_gp5_arcache,
input  wire [2:0]    consumer_axi_gp5_arprot, 
input  wire          consumer_axi_gp5_arvalid,
output wire          consumer_axi_gp5_arready,
output wire [5:0]    consumer_axi_gp5_rid,    
output wire [127:0]  consumer_axi_gp5_rdata,  
output wire [1:0]    consumer_axi_gp5_rresp,  
output wire          consumer_axi_gp5_rlast,  
output wire          consumer_axi_gp5_rvalid, 
input  wire          consumer_axi_gp5_rready, 
input  wire [3:0]    consumer_axi_gp5_awqos,  
input  wire [3:0]    consumer_axi_gp5_arqos,  
output wire [7:0]    consumer_axi_gp5_rcount, 
output wire [7:0]    consumer_axi_gp5_wcount, 
output wire [3:0]    consumer_axi_gp5_racount,
output wire [3:0]    consumer_axi_gp5_wacount,

input  wire          consumer_axi_gp6_aruser,
input  wire          consumer_axi_gp6_awuser, 
input  wire [5:0]    consumer_axi_gp6_awid,   
input  wire [48:0]   consumer_axi_gp6_awaddr, 
input  wire [7:0]    consumer_axi_gp6_awlen , 
input  wire [2:0]    consumer_axi_gp6_awsize, 
input  wire [1:0]    consumer_axi_gp6_awburst,
input  wire          consumer_axi_gp6_awlock, 
input  wire [3:0]    consumer_axi_gp6_awcache,
input  wire [2:0]    consumer_axi_gp6_awprot, 
input  wire          consumer_axi_gp6_awvalid,
output wire          consumer_axi_gp6_awready,
input  wire [127:0]  consumer_axi_gp6_wdata,  
input  wire [15:0]   consumer_axi_gp6_wstrb, 
input  wire          consumer_axi_gp6_wlast,  
input  wire          consumer_axi_gp6_wvalid, 
output wire          consumer_axi_gp6_wready, 
output wire [5:0]    consumer_axi_gp6_bid,    
output wire [1:0]    consumer_axi_gp6_bresp,  
output wire          consumer_axi_gp6_bvalid, 
input  wire          consumer_axi_gp6_bready, 
input  wire [5:0]    consumer_axi_gp6_arid,   
input  wire [48:0]   consumer_axi_gp6_araddr, 
input  wire [7:0]    consumer_axi_gp6_arlen,  
input  wire [2:0]    consumer_axi_gp6_arsize, 
input  wire [1:0]    consumer_axi_gp6_arburst,
input  wire          consumer_axi_gp6_arlock, 
input  wire [3:0]    consumer_axi_gp6_arcache,
input  wire [2:0]    consumer_axi_gp6_arprot, 
input  wire          consumer_axi_gp6_arvalid,
output wire          consumer_axi_gp6_arready,
output wire [5:0]    consumer_axi_gp6_rid,    
output wire [127:0]  consumer_axi_gp6_rdata,  
output wire [1:0]    consumer_axi_gp6_rresp,  
output wire          consumer_axi_gp6_rlast,  
output wire          consumer_axi_gp6_rvalid, 
input  wire          consumer_axi_gp6_rready, 
input  wire [3:0]    consumer_axi_gp6_awqos,  
input  wire [3:0]    consumer_axi_gp6_arqos,  
output wire [7:0]    consumer_axi_gp6_rcount, 
output wire [7:0]    consumer_axi_gp6_wcount, 
output wire [3:0]    consumer_axi_gp6_racount,
output wire [3:0]    consumer_axi_gp6_wacount,

input  wire [39:0]   consumer_axi_acp_awaddr,
input  wire [4:0]    consumer_axi_acp_awid,
input  wire [7:0]    consumer_axi_acp_awlen,
input  wire [2:0]    consumer_axi_acp_awsize,
input  wire [1:0]    consumer_axi_acp_awburst,
input  wire          consumer_axi_acp_awlock,
input  wire [3:0]    consumer_axi_acp_awcache,
input  wire [2:0]    consumer_axi_acp_awprot,
input  wire          consumer_axi_acp_awvalid,
output wire          consumer_axi_acp_awready,
input  wire [1:0]    consumer_axi_acp_awuser,
input  wire [3:0]    consumer_axi_acp_awqos,
input  wire          consumer_axi_acp_wlast,
input  wire [127:0]  consumer_axi_acp_wdata,
input  wire [15:0]   consumer_axi_acp_wstrb,
input  wire          consumer_axi_acp_wvalid,
output wire          consumer_axi_acp_wready,
output wire [1:0]    consumer_axi_acp_bresp,
output wire [4:0]    consumer_axi_acp_bid,
output wire          consumer_axi_acp_bvalid,
input  wire          consumer_axi_acp_bready,
input  wire [39:0]   consumer_axi_acp_araddr,
input  wire [4:0]    consumer_axi_acp_arid,
input  wire [7:0]    consumer_axi_acp_arlen,
input  wire [2:0]    consumer_axi_acp_arsize,
input  wire [1:0]    consumer_axi_acp_arburst,
input  wire          consumer_axi_acp_arlock,
input  wire [3:0]    consumer_axi_acp_arcache,
input  wire [2:0]    consumer_axi_acp_arprot,
input  wire          consumer_axi_acp_arvalid,
output wire          consumer_axi_acp_arready,
input  wire [1:0]    consumer_axi_acp_aruser,
input  wire [3:0]    consumer_axi_acp_arqos,
output wire [4:0]    consumer_axi_acp_rid,
output wire          consumer_axi_acp_rlast,
output wire [127:0]  consumer_axi_acp_rdata,
output wire [1:0]    consumer_axi_acp_rresp,
output wire          consumer_axi_acp_rvalid,
input  wire          consumer_axi_acp_rready,

input  wire [15:0]   consumer_axi_ace_fpd_awuser,
input  wire [15:0]   consumer_axi_ace_fpd_aruser,
input  wire          consumer_axi_ace_fpd_awvalid,
output wire          consumer_axi_ace_fpd_awready,
input  wire [5:0]    consumer_axi_ace_fpd_awid,
input  wire [43:0]   consumer_axi_ace_fpd_awaddr,
input  wire [3:0]    consumer_axi_ace_fpd_awregion,
input  wire [7:0]    consumer_axi_ace_fpd_awlen,
input  wire [2:0]    consumer_axi_ace_fpd_awsize,
input  wire [1:0]    consumer_axi_ace_fpd_awburst,
input  wire          consumer_axi_ace_fpd_awlock,
input  wire [3:0]    consumer_axi_ace_fpd_awcache,
input  wire [2:0]    consumer_axi_ace_fpd_awprot,
input  wire [1:0]    consumer_axi_ace_fpd_awdomain,
input  wire [2:0]    consumer_axi_ace_fpd_awsnoop,
input  wire [1:0]    consumer_axi_ace_fpd_awbar,
input  wire [3:0]    consumer_axi_ace_fpd_awqos,
input  wire          consumer_axi_ace_fpd_wvalid,
output wire          consumer_axi_ace_fpd_wready,
input  wire [127:0]  consumer_axi_ace_fpd_wdata,
input  wire [15:0]   consumer_axi_ace_fpd_wstrb,
input  wire          consumer_axi_ace_fpd_wlast,
input  wire          consumer_axi_ace_fpd_wuser,
output wire          consumer_axi_ace_fpd_bvalid,
input  wire          consumer_axi_ace_fpd_bready,
output wire [5:0]    consumer_axi_ace_fpd_bid,
output wire [1:0]    consumer_axi_ace_fpd_bresp,
output wire          consumer_axi_ace_fpd_buser,
input  wire          consumer_axi_ace_fpd_arvalid,
output wire          consumer_axi_ace_fpd_arready,
input  wire [5:0]    consumer_axi_ace_fpd_arid,
input  wire [43:0]   consumer_axi_ace_fpd_araddr,
input  wire [3:0]    consumer_axi_ace_fpd_arregion,
input  wire [7:0]    consumer_axi_ace_fpd_arlen,
input  wire [2:0]    consumer_axi_ace_fpd_arsize,
input  wire [1:0]    consumer_axi_ace_fpd_arburst,
input  wire          consumer_axi_ace_fpd_arlock,
input  wire [3:0]    consumer_axi_ace_fpd_arcache,
input  wire [2:0]    consumer_axi_ace_fpd_arprot,
input  wire [1:0]    consumer_axi_ace_fpd_ardomain,
input  wire [3:0]    consumer_axi_ace_fpd_arsnoop,
input  wire [1:0]    consumer_axi_ace_fpd_arbar,
input  wire [3:0]    consumer_axi_ace_fpd_arqos,
output wire          consumer_axi_ace_fpd_rvalid,
input  wire          consumer_axi_ace_fpd_rready,
output wire [5:0]    consumer_axi_ace_fpd_rid,
output wire [127:0]  consumer_axi_ace_fpd_rdata,
output wire [3:0]    consumer_axi_ace_fpd_rresp,
output wire          consumer_axi_ace_fpd_rlast,
output wire          consumer_axi_ace_fpd_ruser,
output wire          consumer_axi_ace_fpd_acvalid,
input  wire          consumer_axi_ace_fpd_acready,
output wire [43:0]   consumer_axi_ace_fpd_acaddr,
output wire [3:0]    consumer_axi_ace_fpd_acsnoop,
output wire [2:0]    consumer_axi_ace_fpd_acprot,
input  wire          consumer_axi_ace_fpd_crvalid,
output wire          consumer_axi_ace_fpd_crready,
input  wire [4:0]    consumer_axi_ace_fpd_crresp,
input  wire          consumer_axi_ace_fpd_cdvalid,
output wire          consumer_axi_ace_fpd_cdready,
input  wire [127:0]  consumer_axi_ace_fpd_cddata,
input  wire          consumer_axi_ace_fpd_cdlast,
input  wire          consumer_axi_ace_fpd_wack,
input  wire          consumer_axi_ace_fpd_rack,

// supplier and consumer dp audio axi streams
input  wire [31:0] consumer_axi_stream_dp_audio_tdata,
input  wire consumer_axi_stream_dp_audio_tid,
input  wire consumer_axi_stream_dp_audio_tvalid,
output wire consumer_axi_stream_dp_audio_tready,
output wire [31:0] supplier_axi_stream_dp_mixed_audio_tdata,
output wire supplier_axi_stream_dp_mixed_audio_tid,
output wire supplier_axi_stream_dp_mixed_audio_tvalid,
input  wire supplier_axi_stream_dp_mixed_audio_tready,


// emio ports
output wire emio_can0_phy_tx,
input  wire emio_can0_phy_rx,

output wire emio_can1_phy_tx,
input  wire emio_can1_phy_rx,

output wire [2:0] emio_enet0_speed_mode,
input  wire emio_enet0_gmii_crs,
input  wire emio_enet0_gmii_col,
input  wire [7:0] emio_enet0_gmii_rxd,
input  wire emio_enet0_gmii_rx_er,
input  wire emio_enet0_gmii_rx_dv,
output wire [7:0] emio_enet0_gmii_txd,
output wire emio_enet0_gmii_tx_en,
output wire emio_enet0_gmii_tx_er,
output wire emio_enet0_mdio_mdc,
input  wire emio_enet0_mdio_i,
output wire emio_enet0_mdio_o,
output wire emio_enet0_mdio_t_n,

output wire [2:0] emio_enet1_speed_mode,
input  wire emio_enet1_gmii_crs,
input  wire emio_enet1_gmii_col,
input  wire [7:0] emio_enet1_gmii_rxd,
input  wire emio_enet1_gmii_rx_er,
input  wire emio_enet1_gmii_rx_dv,
output wire [7:0] emio_enet1_gmii_txd,
output wire emio_enet1_gmii_tx_en,
output wire emio_enet1_gmii_tx_er,
output wire emio_enet1_mdio_mdc,
input  wire emio_enet1_mdio_i,
output wire emio_enet1_mdio_o,
output wire emio_enet1_mdio_t_n,

output wire [2:0] emio_enet2_speed_mode,
input  wire emio_enet2_gmii_crs,
input  wire emio_enet2_gmii_col,
input  wire [7:0] emio_enet2_gmii_rxd,
input  wire emio_enet2_gmii_rx_er,
input  wire emio_enet2_gmii_rx_dv,
output wire [7:0] emio_enet2_gmii_txd,
output wire emio_enet2_gmii_tx_en,
output wire emio_enet2_gmii_tx_er,
output wire emio_enet2_mdio_mdc,
input  wire emio_enet2_mdio_i,
output wire emio_enet2_mdio_o,
output wire emio_enet2_mdio_t_n,

output wire [2:0] emio_enet3_speed_mode,
input  wire emio_enet3_gmii_crs,
input  wire emio_enet3_gmii_col,
input  wire [7:0] emio_enet3_gmii_rxd,
output wire [7:0] emio_enet3_gmii_txd,
output wire emio_enet3_gmii_tx_en,
output wire emio_enet3_gmii_tx_er,
output wire emio_enet3_mdio_mdc,
input  wire emio_enet3_mdio_i,
output wire emio_enet3_mdio_o,
output wire emio_enet3_mdio_t_n,

input  wire emio_enet0_tx_r_data_rdy,
output wire emio_enet0_tx_r_rd,
input  wire emio_enet0_tx_r_valid,
input  wire [7:0] emio_enet0_tx_r_data,
input  wire emio_enet0_tx_r_sop,
input  wire emio_enet0_tx_r_eop,
input  wire emio_enet0_tx_r_err,
input  wire emio_enet0_tx_r_underflow,
input  wire emio_enet0_tx_r_flushed,
input  wire emio_enet0_tx_r_control,
output wire emio_enet0_dma_tx_end_tog,
input  wire emio_enet0_dma_tx_status_tog,
output wire [3:0] emio_enet0_tx_r_status,
output wire emio_enet0_rx_w_wr,
output wire [7:0] emio_enet0_rx_w_data,
output wire emio_enet0_rx_w_sop,
output wire emio_enet0_rx_w_eop,
output wire [44:0] emio_enet0_rx_w_status,
output wire emio_enet0_rx_w_err,
input  wire emio_enet0_rx_w_overflow,
input  wire emio_enet0_signal_detect,
output wire emio_enet0_rx_w_flush,
output wire emio_enet0_tx_r_fixed_lat,

input  wire emio_enet1_tx_r_data_rdy,
output wire emio_enet1_tx_r_rd,
input  wire emio_enet1_tx_r_valid,
input  wire [7:0] emio_enet1_tx_r_data,
input  wire emio_enet1_tx_r_sop,
input  wire emio_enet1_tx_r_eop,
input  wire emio_enet1_tx_r_err,
input  wire emio_enet1_tx_r_underflow,
input  wire emio_enet1_tx_r_flushed,
input  wire emio_enet1_tx_r_control,
output wire emio_enet1_dma_tx_end_tog,
input  wire emio_enet1_dma_tx_status_tog,
output wire [3:0] emio_enet1_tx_r_status,
output wire emio_enet1_rx_w_wr,
output wire [7:0] emio_enet1_rx_w_data,
output wire emio_enet1_rx_w_sop,
output wire emio_enet1_rx_w_eop,
output wire [44:0] emio_enet1_rx_w_status,
output wire emio_enet1_rx_w_err,
input  wire emio_enet1_rx_w_overflow,
input  wire emio_enet1_signal_detect,
output wire emio_enet1_rx_w_flush,
output wire emio_enet1_tx_r_fixed_lat,

input  wire emio_enet2_tx_r_data_rdy,
output wire emio_enet2_tx_r_rd,
input  wire emio_enet2_tx_r_valid,
input  wire [7:0] emio_enet2_tx_r_data,
input  wire emio_enet2_tx_r_sop,
input  wire emio_enet2_tx_r_eop,
input  wire emio_enet2_tx_r_err,
input  wire emio_enet2_tx_r_underflow,
input  wire emio_enet2_tx_r_flushed,
input  wire emio_enet2_tx_r_control,
output wire emio_enet2_dma_tx_end_tog,
input  wire emio_enet2_dma_tx_status_tog,
output wire [3:0] emio_enet2_tx_r_status,
output wire emio_enet2_rx_w_wr,
output wire [7:0] emio_enet2_rx_w_data,
output wire emio_enet2_rx_w_sop,
output wire emio_enet2_rx_w_eop,
output wire [44:0] emio_enet2_rx_w_status,
output wire emio_enet2_rx_w_err,
input  wire emio_enet2_rx_w_overflow,
input  wire emio_enet2_signal_detect,
output wire emio_enet2_rx_w_flush,
output wire emio_enet2_tx_r_fixed_lat,

input  wire emio_enet3_tx_r_data_rdy,
output wire emio_enet3_tx_r_rd,
input  wire emio_enet3_tx_r_valid,
input  wire [7:0] emio_enet3_tx_r_data,
input  wire emio_enet3_tx_r_sop,
input  wire emio_enet3_tx_r_eop,
input  wire emio_enet3_tx_r_err,
input  wire emio_enet3_tx_r_underflow,
input  wire emio_enet3_tx_r_flushed,
input  wire emio_enet3_tx_r_control,
output wire emio_enet3_dma_tx_end_tog,
input  wire emio_enet3_dma_tx_status_tog,
output wire [3:0] emio_enet3_tx_r_status,
output wire emio_enet3_rx_w_wr,
output wire [7:0] emio_enet3_rx_w_data,
output wire emio_enet3_rx_w_sop,
output wire emio_enet3_rx_w_eop,
output wire [44:0] emio_enet3_rx_w_status,
output wire emio_enet3_rx_w_err,
input  wire emio_enet3_rx_w_overflow,
input  wire emio_enet3_signal_detect,
output wire emio_enet3_rx_w_flush,
output wire emio_enet3_tx_r_fixed_lat,

output wire emio_enet0_tx_sof,
output wire emio_enet0_sync_frame_tx,
output wire emio_enet0_delay_req_tx,
output wire emio_enet0_pdelay_req_tx,
output wire emio_enet0_pdelay_resp_tx,
output wire emio_enet0_rx_sof,
output wire emio_enet0_sync_frame_rx,
output wire emio_enet0_delay_req_rx,
output wire emio_enet0_pdelay_req_rx,
output wire emio_enet0_pdelay_resp_rx,
input  wire [1:0] emio_enet0_tsu_inc_ctrl,
output wire emio_enet0_tsu_timer_cmp_val,
output wire emio_enet1_tx_sof,
output wire emio_enet1_sync_frame_tx,
output wire emio_enet1_delay_req_tx,
output wire emio_enet1_pdelay_req_tx,
output wire emio_enet1_pdelay_resp_tx,
output wire emio_enet1_rx_sof,
output wire emio_enet1_sync_frame_rx,
output wire emio_enet1_delay_req_rx,
output wire emio_enet1_pdelay_req_rx,
output wire emio_enet1_pdelay_resp_rx,
input  wire [1:0] emio_enet1_tsu_inc_ctrl,
output wire emio_enet1_tsu_timer_cmp_val,
output wire emio_enet2_tx_sof,
output wire emio_enet2_sync_frame_tx,
output wire emio_enet2_delay_req_tx,
output wire emio_enet2_pdelay_req_tx,
output wire emio_enet2_pdelay_resp_tx,
output wire emio_enet2_rx_sof,
output wire emio_enet2_sync_frame_rx,
output wire emio_enet2_delay_req_rx,
output wire emio_enet2_pdelay_req_rx,
output wire emio_enet2_pdelay_resp_rx,
input  wire [1:0] emio_enet2_tsu_inc_ctrl,
output wire emio_enet2_tsu_timer_cmp_val,
output wire emio_enet3_tx_sof,
output wire emio_enet3_sync_frame_tx,
output wire emio_enet3_delay_req_tx,
output wire emio_enet3_pdelay_req_tx,
output wire emio_enet3_pdelay_resp_tx,
output wire emio_enet3_rx_sof,
output wire emio_enet3_sync_frame_rx,
output wire emio_enet3_delay_req_rx,
output wire emio_enet3_pdelay_req_rx,
output wire emio_enet3_pdelay_resp_rx,
input  wire [1:0] emio_enet3_tsu_inc_ctrl,
output wire emio_enet3_tsu_timer_cmp_val,

input  wire emio_enet3_gmii_rx_er,
input  wire emio_enet3_gmii_rx_dv,
output wire [93:0] emio_enet0_enet_tsu_timer_cnt,
input  wire emio_enet0_ext_int_in,
input  wire emio_enet1_ext_int_in,
input  wire emio_enet2_ext_int_in,
input  wire emio_enet3_ext_int_in,
output wire [1:0] emio_enet0_dma_bus_width,
output wire [1:0] emio_enet1_dma_bus_width,
output wire [1:0] emio_enet2_dma_bus_width,
output wire [1:0] emio_enet3_dma_bus_width,

input  wire [95:0] emio_gpio_i,
output wire [95:0] emio_gpio_o,
output wire [95:0] emio_gpio_t_n,

input  wire emio_i2c0_scl_i,
output wire emio_i2c0_scl_o,
output wire emio_i2c0_scl_t_n,
input  wire emio_i2c0_sda_i,
output wire emio_i2c0_sda_o,
output wire emio_i2c0_sda_t_n,

input  wire emio_i2c1_scl_i,
output wire emio_i2c1_scl_o,
output wire emio_i2c1_scl_t_n,
input  wire emio_i2c1_sda_i,
output wire emio_i2c1_sda_o,
output wire emio_i2c1_sda_t_n,

output wire emio_uart0_txd,
input  wire emio_uart0_rxd,
input  wire emio_uart0_ctsn,
output wire emio_uart0_rtsn,
input  wire emio_uart0_dsrn,
input  wire emio_uart0_dcdn,
input  wire emio_uart0_rin,
output wire emio_uart0_dtrn,

output wire emio_uart1_txd,
input  wire emio_uart1_rxd, 
input  wire emio_uart1_ctsn,
output wire emio_uart1_rtsn,
input  wire emio_uart1_dsrn,
input  wire emio_uart1_dcdn,
input  wire emio_uart1_rin, 
output wire emio_uart1_dtrn,

output wire emio_sdio0_cmdout,
input  wire emio_sdio0_cmdin,
output wire emio_sdio0_cmdena_n,
input  wire [7:0] emio_sdio0_datain,
output wire [7:0] emio_sdio0_dataout,
output wire [7:0] emio_sdio0_dataena_n,
input  wire emio_sdio0_cd_n,
input  wire emio_sdio0_wp,
output wire emio_sdio0_ledcontrol,
output wire emio_sdio0_buspower,
output wire [2:0] emio_sdio0_bus_volt,

output wire emio_sdio1_cmdout,        
input  wire emio_sdio1_cmdin,         
output wire emio_sdio1_cmdena_n,        
input  wire [7:0] emio_sdio1_datain,  
output wire [7:0] emio_sdio1_dataout, 
output wire [7:0] emio_sdio1_dataena_n, 
input  wire emio_sdio1_cd_n,          
input  wire emio_sdio1_wp,            
output wire emio_sdio1_ledcontrol,    
output wire emio_sdio1_buspower,      
output wire [2:0] emio_sdio1_bus_volt,

input  wire emio_spi0_m_i,
output wire emio_spi0_m_o,
output wire emio_spi0_mo_t_n,
input  wire emio_spi0_s_i,
output wire emio_spi0_s_o,
output wire emio_spi0_so_t_n,
input  wire emio_spi0_ss_i_n,
output wire emio_spi0_ss_o_n,
output wire emio_spi0_ss1_o_n,
output wire emio_spi0_ss2_o_n,
output wire emio_spi0_ss_n_t_n,
input  wire emio_spi0_sclk_i,
output wire emio_spi0_sclk_o,
output wire emio_spi0_sclk_t_n,
   
input  wire emio_spi1_m_i,         
output wire emio_spi1_m_o,         
output wire emio_spi1_mo_t_n,      
input  wire emio_spi1_s_i,         
output wire emio_spi1_s_o,         
output wire emio_spi1_so_t_n,      
input  wire emio_spi1_ss_i_n,      
output wire emio_spi1_ss_o_n,
output wire emio_spi1_ss1_o_n,
output wire emio_spi1_ss2_o_n,
output wire emio_spi1_ss_n_t_n,    
input  wire emio_spi1_sclk_i,
output wire emio_spi1_sclk_o,      
output wire emio_spi1_sclk_t_n, 

output wire ps_pl_tracectl,
output wire [31:0] ps_pl_tracedata,

output wire [2:0] emio_ttc0_wave_o,
output wire [2:0] emio_ttc1_wave_o,
output wire [2:0] emio_ttc2_wave_o,
output wire [2:0] emio_ttc3_wave_o,

output wire emio_wdt0_rst_o,
output wire emio_wdt1_rst_o,

input  wire emio_hub_port_overcrnt_usb3_0,
input  wire emio_hub_port_overcrnt_usb3_1,
input  wire emio_hub_port_overcrnt_usb2_0,
input  wire emio_hub_port_overcrnt_usb2_1,
output wire emio_u2dsport_vbus_ctrl_usb3_0,
output wire emio_u2dsport_vbus_ctrl_usb3_1,
output wire emio_u3dsport_vbus_ctrl_usb3_0,
output wire emio_u3dsport_vbus_ctrl_usb3_1,

input  wire [7:0] pl2adma_cvld,
input  wire [7:0] pl2adma_tack,
output wire [7:0] adma2pl_cack,
output wire [7:0] adma2pl_tvld,

input  wire [7:0] perif_gdma_cvld,
input  wire [7:0] perif_gdma_tack,
output wire [7:0] gdma_perif_cack,
output wire [7:0] gdma_perif_tvld,

input  wire [3:0] pl_clock_stop,

input  wire dp_live_video_in_vsync,
input  wire dp_live_video_in_hsync,
input  wire dp_live_video_in_de,
input  wire [35:0] dp_live_video_in_pixel1,
output wire dp_video_out_hsync,
output wire dp_video_out_vsync,
output wire [35:0] dp_video_out_pixel1,
input  wire dp_aux_data_in,
output wire dp_aux_data_out,
output wire dp_aux_data_oe_n,
input  wire [7:0] dp_live_gfx_alpha_in,
input  wire [35:0] dp_live_gfx_pixel1_in,
input  wire dp_hot_plug_detect,
input  wire dp_external_custom_event1,
input  wire dp_external_custom_event2,
input  wire dp_external_vsync_event,
output wire dp_live_video_de_out, 	

input  wire pl_ps_eventi,
output wire ps_pl_evento,
output wire [3:0] ps_pl_standbywfe,
output wire [3:0] ps_pl_standbywfi,
input  wire [3:0] pl_ps_apugic_irq,
input  wire [3:0] pl_ps_apugic_fiq,

input  wire rpu_eventi0,
input  wire rpu_eventi1,
output wire rpu_evento0,
output wire rpu_evento1,
input  wire nfiq0_lpd_rpu,
input  wire nfiq1_lpd_rpu,
input  wire nirq0_lpd_rpu,
input  wire nirq1_lpd_rpu,

output wire irq_ipi_pl_0,
output wire irq_ipi_pl_1,
output wire irq_ipi_pl_2,
output wire irq_ipi_pl_3,

input  wire [59:0] stm_event,

// ftm
input  wire [3:0] pl_ps_trigack,
input  wire [3:0] pl_ps_trigger,
output wire [3:0] ps_pl_trigack,
output wire [3:0] ps_pl_trigger,
output wire [31:0] ftm_gpo,
input  wire [31:0] ftm_gpi,

input  wire [7:0] pl_ps_irq0,
input  wire [7:0] pl_ps_irq1,

output wire fps_tpl_reset0_n,
output wire fps_tpl_reset1_n,
output wire fps_tpl_reset2_n,
output wire fps_tpl_reset3_n,

output wire fps_tpl_irq_can0,
output wire fps_tpl_irq_can1,
output wire fps_tpl_irq_enet0,
output wire fps_tpl_irq_enet1,
output wire fps_tpl_irq_enet2,
output wire fps_tpl_irq_enet3,
output wire fps_tpl_irq_enet0_wake,
output wire fps_tpl_irq_enet1_wake,
output wire fps_tpl_irq_enet2_wake,
output wire fps_tpl_irq_enet3_wake,
output wire fps_tpl_irq_gpio,
output wire fps_tpl_irq_i2c0,
output wire fps_tpl_irq_i2c1,
output wire fps_tpl_irq_uart0,
output wire fps_tpl_irq_uart1,
output wire fps_tpl_irq_sdio0,
output wire fps_tpl_irq_sdio1,
output wire fps_tpl_irq_sdio0_wake,
output wire fps_tpl_irq_sdio1_wake,
output wire fps_tpl_irq_spi0,
output wire fps_tpl_irq_spi1,
output wire fps_tpl_irq_qspi,
output wire fps_tpl_irq_ttc0_0,
output wire fps_tpl_irq_ttc0_1,
output wire fps_tpl_irq_ttc0_2,
output wire fps_tpl_irq_ttc1_0,
output wire fps_tpl_irq_ttc1_1,
output wire fps_tpl_irq_ttc1_2,
output wire fps_tpl_irq_ttc2_0,
output wire fps_tpl_irq_ttc2_1,
output wire fps_tpl_irq_ttc2_2,
output wire fps_tpl_irq_ttc3_0,
output wire fps_tpl_irq_ttc3_1,
output wire fps_tpl_irq_ttc3_2,
output wire fps_tpl_irq_csu_pmu_wdt,
output wire fps_tpl_irq_lp_wdt,
output wire [3:0] fps_tpl_irq_usb3_0_endpoint,
output wire fps_tpl_irq_usb3_0_otg,
output wire [3:0] fps_tpl_irq_usb3_1_endpoint,
output wire fps_tpl_irq_usb3_1_otg,
output wire [7:0] fps_tpl_irq_adma_chan,
output wire [1:0] fps_tpl_irq_usb3_0_pmu_wakeup,
output wire [7:0] fps_tpl_irq_gdma_chan,
output wire fps_tpl_irq_csu,
output wire fps_tpl_irq_csu_dma,
output wire fps_tpl_irq_efuse,
output wire fps_tpl_irq_xmpu_lpd,
output wire fps_tpl_irq_ddr_ss,
output wire fps_tpl_irq_nand,
output wire fps_tpl_irq_fp_wdt,
output wire [1:0] fps_tpl_irq_pcie_msi, 
output wire fps_tpl_irq_pcie_legacy, 
output wire fps_tpl_irq_pcie_dma, 
output wire fps_tpl_irq_pcie_msc, 
output wire fps_tpl_irq_dport, 
output wire fps_tpl_irq_fpd_apb_int, 
output wire fps_tpl_irq_fpd_atb_error, 
output wire fps_tpl_irq_dpdma, 
output wire fps_tpl_irq_apm_fpd, 
output wire fps_tpl_irq_gpu, 
output wire fps_tpl_irq_sata, 
output wire fps_tpl_irq_xmpu_fpd, 
output wire [3:0] fps_tpl_irq_apu_cpumnt, 
output wire [3:0] fps_tpl_irq_apu_cti, 
output wire [3:0] fps_tpl_irq_apu_pmu, 
output wire [3:0] fps_tpl_irq_apu_comm, 
output wire fps_tpl_irq_apu_l2err, 
output wire fps_tpl_irq_apu_exterr, 
output wire fps_tpl_irq_apu_regs, 
output wire fps_tpl_irq_intf_ppd_cci, 
output wire fps_tpl_irq_intf_fpd_smmu,
output wire fps_tpl_irq_atb_err_lpd,
output wire fps_tpl_irq_aib_axi,
output wire fps_tpl_irq_ams,
output wire fps_tpl_irq_lpd_apm,
output wire fps_tpl_irq_rtc_alaram,
output wire fps_tpl_irq_rtc_seconds,
output wire fps_tpl_irq_clkmon,
output wire fps_tpl_irq_ipi_channel0,
output wire fps_tpl_irq_ipi_channel1,
output wire fps_tpl_irq_ipi_channel2,
output wire fps_tpl_irq_ipi_channel7,
output wire fps_tpl_irq_ipi_channel8,
output wire fps_tpl_irq_ipi_channel9,
output wire fps_tpl_irq_ipi_channel10,
output wire [1:0] fps_tpl_irq_rpu_pm,
output wire fps_tpl_irq_ocm_error,
output wire fps_tpl_irq_lpd_apb_intr,
output wire fps_tpl_irq_r5_core0_ecc_error,
output wire fps_tpl_irq_r5_core1_ecc_error,


output wire osc_rtc_clk,

input  wire [31:0] pl_pmu_gpi,
output wire [31:0] pmu_pl_gpo,
input  wire aib_pmu_afifm_fpd_ack,
input  wire aib_pmu_afifm_lpd_ack,
output wire pmu_aib_afifm_fpd_req,
output wire pmu_aib_afifm_lpd_req,
output wire [46:0] pmu_error_to_pl,
input  wire [3:0] pmu_error_from_pl,

input  wire ddrc_ext_refresh_rank0_req,
input  wire ddrc_ext_refresh_rank1_req,
input  wire pl_acpinact,

input  [31:0] pstp_pl_in,
output [31:0] pstp_pl_out,
input  [31:0] pstp_pl_ts
);

// these are not used sinks for irq lines form PS
wire [18:0] irq_lpd_dev_null;
wire [19:0] irq_fpd_dev_null;

// unclear what these are
wire pss_alto_core_pad_mgttxn0out;
wire pss_alto_core_pad_mgttxp0out;
wire pss_alto_core_pad_mgttxn1out;
wire pss_alto_core_pad_mgttxp1out;
wire pss_alto_core_pad_mgttxn2out;
wire pss_alto_core_pad_mgttxp2out;
wire pss_alto_core_pad_mgttxn3out;
wire pss_alto_core_pad_mgttxp3out;
wire pss_alto_core_pad_pado;

// rename the gpio reset lins
assign fps_tpl_reset0_n = emio_gpio_i[95];
assign fps_tpl_reset1_n = emio_gpio_i[94];
assign fps_tpl_reset2_n = emio_gpio_i[93];
assign fps_tpl_reset3_n = emio_gpio_i[92];

PS8 PS8_i  (
.MAXIGP0ACLK (clk_tps_fpl_supplier_axi_hpm0_fpd),
.MAXIGP0AWID (supplier_axi_gp0_awid),
.MAXIGP0AWADDR (supplier_axi_gp0_awaddr),
.MAXIGP0AWLEN (supplier_axi_gp0_awlen),
.MAXIGP0AWSIZE (supplier_axi_gp0_awsize),
.MAXIGP0AWBURST (supplier_axi_gp0_awburst),
.MAXIGP0AWLOCK (supplier_axi_gp0_awlock),
.MAXIGP0AWCACHE (supplier_axi_gp0_awcache),
.MAXIGP0AWPROT (supplier_axi_gp0_awprot),
.MAXIGP0AWVALID (supplier_axi_gp0_awvalid),
.MAXIGP0AWUSER (supplier_axi_gp0_awuser),
.MAXIGP0AWREADY (supplier_axi_gp0_awready),
.MAXIGP0WDATA (supplier_axi_gp0_wdata),
.MAXIGP0WSTRB (supplier_axi_gp0_wstrb),
.MAXIGP0WLAST (supplier_axi_gp0_wlast),
.MAXIGP0WVALID (supplier_axi_gp0_wvalid),
.MAXIGP0WREADY (supplier_axi_gp0_wready),
.MAXIGP0BID (supplier_axi_gp0_bid),
.MAXIGP0BRESP (supplier_axi_gp0_bresp),
.MAXIGP0BVALID (supplier_axi_gp0_bvalid),
.MAXIGP0BREADY (supplier_axi_gp0_bready),
.MAXIGP0ARID (supplier_axi_gp0_arid),
.MAXIGP0ARADDR (supplier_axi_gp0_araddr),
.MAXIGP0ARLEN (supplier_axi_gp0_arlen),
.MAXIGP0ARSIZE (supplier_axi_gp0_arsize),
.MAXIGP0ARBURST (supplier_axi_gp0_arburst),
.MAXIGP0ARLOCK (supplier_axi_gp0_arlock),
.MAXIGP0ARCACHE (supplier_axi_gp0_arcache),
.MAXIGP0ARPROT (supplier_axi_gp0_arprot),
.MAXIGP0ARVALID (supplier_axi_gp0_arvalid),
.MAXIGP0ARUSER (supplier_axi_gp0_aruser),
.MAXIGP0ARREADY (supplier_axi_gp0_arready),
.MAXIGP0RID (supplier_axi_gp0_rid),
.MAXIGP0RDATA (supplier_axi_gp0_rdata),
.MAXIGP0RRESP (supplier_axi_gp0_rresp),
.MAXIGP0RLAST (supplier_axi_gp0_rlast),
.MAXIGP0RVALID (supplier_axi_gp0_rvalid),
.MAXIGP0RREADY (supplier_axi_gp0_rready),
.MAXIGP0AWQOS (supplier_axi_gp0_awqos),
.MAXIGP0ARQOS (supplier_axi_gp0_arqos),
.MAXIGP1ACLK (clk_tps_fpl_supplier_axi_hpm1_fpd),
.MAXIGP1AWID (supplier_axi_gp1_awid),
.MAXIGP1AWADDR (supplier_axi_gp1_awaddr),
.MAXIGP1AWLEN (supplier_axi_gp1_awlen),
.MAXIGP1AWSIZE (supplier_axi_gp1_awsize),
.MAXIGP1AWBURST (supplier_axi_gp1_awburst),
.MAXIGP1AWLOCK (supplier_axi_gp1_awlock),
.MAXIGP1AWCACHE (supplier_axi_gp1_awcache),
.MAXIGP1AWPROT (supplier_axi_gp1_awprot),
.MAXIGP1AWVALID (supplier_axi_gp1_awvalid),
.MAXIGP1AWUSER (supplier_axi_gp1_awuser),
.MAXIGP1AWREADY (supplier_axi_gp1_awready),
.MAXIGP1WDATA (supplier_axi_gp1_wdata),
.MAXIGP1WSTRB (supplier_axi_gp1_wstrb),
.MAXIGP1WLAST (supplier_axi_gp1_wlast),
.MAXIGP1WVALID (supplier_axi_gp1_wvalid),
.MAXIGP1WREADY (supplier_axi_gp1_wready),
.MAXIGP1BID (supplier_axi_gp1_bid),
.MAXIGP1BRESP (supplier_axi_gp1_bresp),
.MAXIGP1BVALID (supplier_axi_gp1_bvalid),
.MAXIGP1BREADY (supplier_axi_gp1_bready),
.MAXIGP1ARID (supplier_axi_gp1_arid),
.MAXIGP1ARADDR (supplier_axi_gp1_araddr),
.MAXIGP1ARLEN (supplier_axi_gp1_arlen),
.MAXIGP1ARSIZE (supplier_axi_gp1_arsize),
.MAXIGP1ARBURST (supplier_axi_gp1_arburst),
.MAXIGP1ARLOCK (supplier_axi_gp1_arlock),
.MAXIGP1ARCACHE (supplier_axi_gp1_arcache),
.MAXIGP1ARPROT (supplier_axi_gp1_arprot),
.MAXIGP1ARVALID (supplier_axi_gp1_arvalid),
.MAXIGP1ARUSER (supplier_axi_gp1_aruser),
.MAXIGP1ARREADY (supplier_axi_gp1_arready),
.MAXIGP1RID (supplier_axi_gp1_rid),
.MAXIGP1RDATA (supplier_axi_gp1_rdata),
.MAXIGP1RRESP (supplier_axi_gp1_rresp),
.MAXIGP1RLAST (supplier_axi_gp1_rlast),
.MAXIGP1RVALID (supplier_axi_gp1_rvalid),
.MAXIGP1RREADY (supplier_axi_gp1_rready),
.MAXIGP1AWQOS (supplier_axi_gp1_awqos),
.MAXIGP1ARQOS (supplier_axi_gp1_arqos),
.MAXIGP2ACLK (clk_tps_fpl_supplier_axi_hpm0_lpd),
.MAXIGP2AWID (supplier_axi_gp2_awid),
.MAXIGP2AWADDR (supplier_axi_gp2_awaddr),
.MAXIGP2AWLEN (supplier_axi_gp2_awlen),
.MAXIGP2AWSIZE (supplier_axi_gp2_awsize),
.MAXIGP2AWBURST (supplier_axi_gp2_awburst),
.MAXIGP2AWLOCK (supplier_axi_gp2_awlock),
.MAXIGP2AWCACHE (supplier_axi_gp2_awcache),
.MAXIGP2AWPROT (supplier_axi_gp2_awprot),
.MAXIGP2AWVALID (supplier_axi_gp2_awvalid),
.MAXIGP2AWUSER (supplier_axi_gp2_awuser),
.MAXIGP2AWREADY (supplier_axi_gp2_awready),
.MAXIGP2WDATA (supplier_axi_gp2_wdata),
.MAXIGP2WSTRB (supplier_axi_gp2_wstrb),
.MAXIGP2WLAST (supplier_axi_gp2_wlast),
.MAXIGP2WVALID (supplier_axi_gp2_wvalid),
.MAXIGP2WREADY (supplier_axi_gp2_wready),
.MAXIGP2BID (supplier_axi_gp2_bid),
.MAXIGP2BRESP (supplier_axi_gp2_bresp),
.MAXIGP2BVALID (supplier_axi_gp2_bvalid),
.MAXIGP2BREADY (supplier_axi_gp2_bready),
.MAXIGP2ARID (supplier_axi_gp2_arid),
.MAXIGP2ARADDR (supplier_axi_gp2_araddr),
.MAXIGP2ARLEN (supplier_axi_gp2_arlen),
.MAXIGP2ARSIZE (supplier_axi_gp2_arsize),
.MAXIGP2ARBURST (supplier_axi_gp2_arburst),
.MAXIGP2ARLOCK (supplier_axi_gp2_arlock),
.MAXIGP2ARCACHE (supplier_axi_gp2_arcache),
.MAXIGP2ARPROT (supplier_axi_gp2_arprot),
.MAXIGP2ARVALID (supplier_axi_gp2_arvalid),
.MAXIGP2ARUSER (supplier_axi_gp2_aruser),
.MAXIGP2ARREADY (supplier_axi_gp2_arready),
.MAXIGP2RID (supplier_axi_gp2_rid),
.MAXIGP2RDATA (supplier_axi_gp2_rdata),
.MAXIGP2RRESP (supplier_axi_gp2_rresp),
.MAXIGP2RLAST (supplier_axi_gp2_rlast),
.MAXIGP2RVALID (supplier_axi_gp2_rvalid),
.MAXIGP2RREADY (supplier_axi_gp2_rready),
.MAXIGP2AWQOS (supplier_axi_gp2_awqos),
.MAXIGP2ARQOS (supplier_axi_gp2_arqos),
.SAXIGP0RCLK (clk_tps_fpl_consumer_axi_hpc0_fpd_read),
.SAXIGP0WCLK (clk_tps_fpl_consumer_axi_hpc0_fpd_write),
.SAXIGP0ARUSER (consumer_axi_gp0_aruser),
.SAXIGP0AWUSER (consumer_axi_gp0_awuser),
.SAXIGP0AWID (consumer_axi_gp0_awid),
.SAXIGP0AWADDR (consumer_axi_gp0_awaddr),
.SAXIGP0AWLEN (consumer_axi_gp0_awlen),
.SAXIGP0AWSIZE (consumer_axi_gp0_awsize),
.SAXIGP0AWBURST (consumer_axi_gp0_awburst),
.SAXIGP0AWLOCK (consumer_axi_gp0_awlock),
.SAXIGP0AWCACHE (consumer_axi_gp0_awcache),
.SAXIGP0AWPROT (consumer_axi_gp0_awprot),
.SAXIGP0AWVALID (consumer_axi_gp0_awvalid),
.SAXIGP0AWREADY (consumer_axi_gp0_awready),
.SAXIGP0WDATA (consumer_axi_gp0_wdata),
.SAXIGP0WSTRB (consumer_axi_gp0_wstrb),
.SAXIGP0WLAST (consumer_axi_gp0_wlast),
.SAXIGP0WVALID (consumer_axi_gp0_wvalid),
.SAXIGP0WREADY (consumer_axi_gp0_wready),
.SAXIGP0BID (consumer_axi_gp0_bid),
.SAXIGP0BRESP (consumer_axi_gp0_bresp),
.SAXIGP0BVALID (consumer_axi_gp0_bvalid),
.SAXIGP0BREADY (consumer_axi_gp0_bready),
.SAXIGP0ARID (consumer_axi_gp0_arid),
.SAXIGP0ARADDR (consumer_axi_gp0_araddr),
.SAXIGP0ARLEN (consumer_axi_gp0_arlen),
.SAXIGP0ARSIZE (consumer_axi_gp0_arsize),
.SAXIGP0ARBURST (consumer_axi_gp0_arburst),
.SAXIGP0ARLOCK (consumer_axi_gp0_arlock),
.SAXIGP0ARCACHE (consumer_axi_gp0_arcache),
.SAXIGP0ARPROT (consumer_axi_gp0_arprot),
.SAXIGP0ARVALID (consumer_axi_gp0_arvalid),
.SAXIGP0ARREADY (consumer_axi_gp0_arready),
.SAXIGP0RID (consumer_axi_gp0_rid),
.SAXIGP0RDATA (consumer_axi_gp0_rdata),
.SAXIGP0RRESP (consumer_axi_gp0_rresp),
.SAXIGP0RLAST (consumer_axi_gp0_rlast),
.SAXIGP0RVALID (consumer_axi_gp0_rvalid),
.SAXIGP0RREADY (consumer_axi_gp0_rready),
.SAXIGP0AWQOS (consumer_axi_gp0_awqos),
.SAXIGP0ARQOS (consumer_axi_gp0_arqos),
.SAXIGP0RCOUNT (consumer_axi_gp0_rcount),
.SAXIGP0WCOUNT (consumer_axi_gp0_wcount),
.SAXIGP0RACOUNT (consumer_axi_gp0_racount),
.SAXIGP0WACOUNT (consumer_axi_gp0_wacount),
.SAXIGP1RCLK (clk_tps_fpl_consumer_axi_hpc1_fpd_read),
.SAXIGP1WCLK (clk_tps_fpl_consumer_axi_hpc1_fpd_write),
.SAXIGP1ARUSER (consumer_axi_gp1_aruser),
.SAXIGP1AWUSER (consumer_axi_gp1_awuser),
.SAXIGP1AWID (consumer_axi_gp1_awid),
.SAXIGP1AWADDR (consumer_axi_gp1_awaddr),
.SAXIGP1AWLEN (consumer_axi_gp1_awlen),
.SAXIGP1AWSIZE (consumer_axi_gp1_awsize),
.SAXIGP1AWBURST (consumer_axi_gp1_awburst),
.SAXIGP1AWLOCK (consumer_axi_gp1_awlock),
.SAXIGP1AWCACHE (consumer_axi_gp1_awcache),
.SAXIGP1AWPROT (consumer_axi_gp1_awprot),
.SAXIGP1AWVALID (consumer_axi_gp1_awvalid),
.SAXIGP1AWREADY (consumer_axi_gp1_awready),
.SAXIGP1WDATA (consumer_axi_gp1_wdata),
.SAXIGP1WSTRB (consumer_axi_gp1_wstrb),
.SAXIGP1WLAST (consumer_axi_gp1_wlast),
.SAXIGP1WVALID (consumer_axi_gp1_wvalid),
.SAXIGP1WREADY (consumer_axi_gp1_wready),
.SAXIGP1BID (consumer_axi_gp1_bid),
.SAXIGP1BRESP (consumer_axi_gp1_bresp),
.SAXIGP1BVALID (consumer_axi_gp1_bvalid),
.SAXIGP1BREADY (consumer_axi_gp1_bready),
.SAXIGP1ARID (consumer_axi_gp1_arid),
.SAXIGP1ARADDR (consumer_axi_gp1_araddr),
.SAXIGP1ARLEN (consumer_axi_gp1_arlen),
.SAXIGP1ARSIZE (consumer_axi_gp1_arsize),
.SAXIGP1ARBURST (consumer_axi_gp1_arburst),
.SAXIGP1ARLOCK (consumer_axi_gp1_arlock),
.SAXIGP1ARCACHE (consumer_axi_gp1_arcache),
.SAXIGP1ARPROT (consumer_axi_gp1_arprot),
.SAXIGP1ARVALID (consumer_axi_gp1_arvalid),
.SAXIGP1ARREADY (consumer_axi_gp1_arready),
.SAXIGP1RID (consumer_axi_gp1_rid),
.SAXIGP1RDATA (consumer_axi_gp1_rdata),
.SAXIGP1RRESP (consumer_axi_gp1_rresp),
.SAXIGP1RLAST (consumer_axi_gp1_rlast),
.SAXIGP1RVALID (consumer_axi_gp1_rvalid),
.SAXIGP1RREADY (consumer_axi_gp1_rready),
.SAXIGP1AWQOS (consumer_axi_gp1_awqos),
.SAXIGP1ARQOS (consumer_axi_gp1_arqos),
.SAXIGP1RCOUNT (consumer_axi_gp1_rcount),
.SAXIGP1WCOUNT (consumer_axi_gp1_wcount),
.SAXIGP1RACOUNT (consumer_axi_gp1_racount),
.SAXIGP1WACOUNT (consumer_axi_gp1_wacount),
.SAXIGP2RCLK (clk_tps_fpl_consumer_axi_hp0_fpd_read),
.SAXIGP2WCLK (clk_tps_fpl_consumer_axi_hp0_fpd_write),
.SAXIGP2ARUSER (consumer_axi_gp2_aruser),
.SAXIGP2AWUSER (consumer_axi_gp2_awuser),
.SAXIGP2AWID (consumer_axi_gp2_awid),
.SAXIGP2AWADDR (consumer_axi_gp2_awaddr),
.SAXIGP2AWLEN (consumer_axi_gp2_awlen),
.SAXIGP2AWSIZE (consumer_axi_gp2_awsize),
.SAXIGP2AWBURST (consumer_axi_gp2_awburst),
.SAXIGP2AWLOCK (consumer_axi_gp2_awlock),
.SAXIGP2AWCACHE (consumer_axi_gp2_awcache),
.SAXIGP2AWPROT (consumer_axi_gp2_awprot),
.SAXIGP2AWVALID (consumer_axi_gp2_awvalid),
.SAXIGP2AWREADY (consumer_axi_gp2_awready),
.SAXIGP2WDATA (consumer_axi_gp2_wdata),
.SAXIGP2WSTRB (consumer_axi_gp2_wstrb),
.SAXIGP2WLAST (consumer_axi_gp2_wlast),
.SAXIGP2WVALID (consumer_axi_gp2_wvalid),
.SAXIGP2WREADY (consumer_axi_gp2_wready),
.SAXIGP2BID (consumer_axi_gp2_bid),
.SAXIGP2BRESP (consumer_axi_gp2_bresp),
.SAXIGP2BVALID (consumer_axi_gp2_bvalid),
.SAXIGP2BREADY (consumer_axi_gp2_bready),
.SAXIGP2ARID (consumer_axi_gp2_arid),
.SAXIGP2ARADDR (consumer_axi_gp2_araddr),
.SAXIGP2ARLEN (consumer_axi_gp2_arlen),
.SAXIGP2ARSIZE (consumer_axi_gp2_arsize),
.SAXIGP2ARBURST (consumer_axi_gp2_arburst),
.SAXIGP2ARLOCK (consumer_axi_gp2_arlock),
.SAXIGP2ARCACHE (consumer_axi_gp2_arcache),
.SAXIGP2ARPROT (consumer_axi_gp2_arprot),
.SAXIGP2ARVALID (consumer_axi_gp2_arvalid),
.SAXIGP2ARREADY (consumer_axi_gp2_arready),
.SAXIGP2RID (consumer_axi_gp2_rid),
.SAXIGP2RDATA (consumer_axi_gp2_rdata),
.SAXIGP2RRESP (consumer_axi_gp2_rresp),
.SAXIGP2RLAST (consumer_axi_gp2_rlast),
.SAXIGP2RVALID (consumer_axi_gp2_rvalid),
.SAXIGP2RREADY (consumer_axi_gp2_rready),
.SAXIGP2AWQOS (consumer_axi_gp2_awqos),
.SAXIGP2ARQOS (consumer_axi_gp2_arqos),
.SAXIGP2RCOUNT (consumer_axi_gp2_rcount),
.SAXIGP2WCOUNT (consumer_axi_gp2_wcount),
.SAXIGP2RACOUNT (consumer_axi_gp2_racount),
.SAXIGP2WACOUNT (consumer_axi_gp2_wacount),
.SAXIGP3RCLK (clk_tps_fpl_consumer_axi_hp1_fpd_read),
.SAXIGP3WCLK (clk_tps_fpl_consumer_axi_hp1_fpd_write),
.SAXIGP3ARUSER (consumer_axi_gp3_aruser),
.SAXIGP3AWUSER (consumer_axi_gp3_awuser),
.SAXIGP3AWID (consumer_axi_gp3_awid),
.SAXIGP3AWADDR (consumer_axi_gp3_awaddr),
.SAXIGP3AWLEN (consumer_axi_gp3_awlen),
.SAXIGP3AWSIZE (consumer_axi_gp3_awsize),
.SAXIGP3AWBURST (consumer_axi_gp3_awburst),
.SAXIGP3AWLOCK (consumer_axi_gp3_awlock),
.SAXIGP3AWCACHE (consumer_axi_gp3_awcache),
.SAXIGP3AWPROT (consumer_axi_gp3_awprot),
.SAXIGP3AWVALID (consumer_axi_gp3_awvalid),
.SAXIGP3AWREADY (consumer_axi_gp3_awready),
.SAXIGP3WDATA (consumer_axi_gp3_wdata),
.SAXIGP3WSTRB (consumer_axi_gp3_wstrb),
.SAXIGP3WLAST (consumer_axi_gp3_wlast),
.SAXIGP3WVALID (consumer_axi_gp3_wvalid),
.SAXIGP3WREADY (consumer_axi_gp3_wready),
.SAXIGP3BID (consumer_axi_gp3_bid),
.SAXIGP3BRESP (consumer_axi_gp3_bresp),
.SAXIGP3BVALID (consumer_axi_gp3_bvalid),
.SAXIGP3BREADY (consumer_axi_gp3_bready),
.SAXIGP3ARID (consumer_axi_gp3_arid),
.SAXIGP3ARADDR (consumer_axi_gp3_araddr),
.SAXIGP3ARLEN (consumer_axi_gp3_arlen),
.SAXIGP3ARSIZE (consumer_axi_gp3_arsize),
.SAXIGP3ARBURST (consumer_axi_gp3_arburst),
.SAXIGP3ARLOCK (consumer_axi_gp3_arlock),
.SAXIGP3ARCACHE (consumer_axi_gp3_arcache),
.SAXIGP3ARPROT (consumer_axi_gp3_arprot),
.SAXIGP3ARVALID (consumer_axi_gp3_arvalid),
.SAXIGP3ARREADY (consumer_axi_gp3_arready),
.SAXIGP3RID (consumer_axi_gp3_rid),
.SAXIGP3RDATA (consumer_axi_gp3_rdata),
.SAXIGP3RRESP (consumer_axi_gp3_rresp),
.SAXIGP3RLAST (consumer_axi_gp3_rlast),
.SAXIGP3RVALID (consumer_axi_gp3_rvalid),
.SAXIGP3RREADY (consumer_axi_gp3_rready),
.SAXIGP3AWQOS (consumer_axi_gp3_awqos),
.SAXIGP3ARQOS (consumer_axi_gp3_arqos),
.SAXIGP3RCOUNT (consumer_axi_gp3_rcount),
.SAXIGP3WCOUNT (consumer_axi_gp3_wcount),
.SAXIGP3RACOUNT (consumer_axi_gp3_racount),
.SAXIGP3WACOUNT (consumer_axi_gp3_wacount),
.SAXIGP4RCLK (clk_tps_fpl_consumer_axi_hp2_fpd_read),
.SAXIGP4WCLK (clk_tps_fpl_consumer_axi_hp2_fpd_write),
.SAXIGP4ARUSER (consumer_axi_gp4_aruser),
.SAXIGP4AWUSER (consumer_axi_gp4_awuser),
.SAXIGP4AWID (consumer_axi_gp4_awid),
.SAXIGP4AWADDR (consumer_axi_gp4_awaddr),
.SAXIGP4AWLEN (consumer_axi_gp4_awlen),
.SAXIGP4AWSIZE (consumer_axi_gp4_awsize),
.SAXIGP4AWBURST (consumer_axi_gp4_awburst),
.SAXIGP4AWLOCK (consumer_axi_gp4_awlock),
.SAXIGP4AWCACHE (consumer_axi_gp4_awcache),
.SAXIGP4AWPROT (consumer_axi_gp4_awprot),
.SAXIGP4AWVALID (consumer_axi_gp4_awvalid),
.SAXIGP4AWREADY (consumer_axi_gp4_awready),
.SAXIGP4WDATA (consumer_axi_gp4_wdata),
.SAXIGP4WSTRB (consumer_axi_gp4_wstrb),
.SAXIGP4WLAST (consumer_axi_gp4_wlast),
.SAXIGP4WVALID (consumer_axi_gp4_wvalid),
.SAXIGP4WREADY (consumer_axi_gp4_wready),
.SAXIGP4BID (consumer_axi_gp4_bid),
.SAXIGP4BRESP (consumer_axi_gp4_bresp),
.SAXIGP4BVALID (consumer_axi_gp4_bvalid),
.SAXIGP4BREADY (consumer_axi_gp4_bready),
.SAXIGP4ARID (consumer_axi_gp4_arid),
.SAXIGP4ARADDR (consumer_axi_gp4_araddr),
.SAXIGP4ARLEN (consumer_axi_gp4_arlen),
.SAXIGP4ARSIZE (consumer_axi_gp4_arsize),
.SAXIGP4ARBURST (consumer_axi_gp4_arburst),
.SAXIGP4ARLOCK (consumer_axi_gp4_arlock),
.SAXIGP4ARCACHE (consumer_axi_gp4_arcache),
.SAXIGP4ARPROT (consumer_axi_gp4_arprot),
.SAXIGP4ARVALID (consumer_axi_gp4_arvalid),
.SAXIGP4ARREADY (consumer_axi_gp4_arready),
.SAXIGP4RID (consumer_axi_gp4_rid),
.SAXIGP4RDATA (consumer_axi_gp4_rdata),
.SAXIGP4RRESP (consumer_axi_gp4_rresp),
.SAXIGP4RLAST (consumer_axi_gp4_rlast),
.SAXIGP4RVALID (consumer_axi_gp4_rvalid),
.SAXIGP4RREADY (consumer_axi_gp4_rready),
.SAXIGP4AWQOS (consumer_axi_gp4_awqos),
.SAXIGP4ARQOS (consumer_axi_gp4_arqos),
.SAXIGP4RCOUNT (consumer_axi_gp4_rcount),
.SAXIGP4WCOUNT (consumer_axi_gp4_wcount),
.SAXIGP4RACOUNT (consumer_axi_gp4_racount),
.SAXIGP4WACOUNT (consumer_axi_gp4_wacount),
.SAXIGP5RCLK (clk_tps_fpl_consumer_axi_hp3_fpd_read),
.SAXIGP5WCLK (clk_tps_fpl_consumer_axi_hp3_fpd_write),
.SAXIGP5ARUSER (consumer_axi_gp5_aruser),
.SAXIGP5AWUSER (consumer_axi_gp5_awuser),
.SAXIGP5AWID (consumer_axi_gp5_awid),
.SAXIGP5AWADDR (consumer_axi_gp5_awaddr),
.SAXIGP5AWLEN (consumer_axi_gp5_awlen),
.SAXIGP5AWSIZE (consumer_axi_gp5_awsize),
.SAXIGP5AWBURST (consumer_axi_gp5_awburst),
.SAXIGP5AWLOCK (consumer_axi_gp5_awlock),
.SAXIGP5AWCACHE (consumer_axi_gp5_awcache),
.SAXIGP5AWPROT (consumer_axi_gp5_awprot),
.SAXIGP5AWVALID (consumer_axi_gp5_awvalid),
.SAXIGP5AWREADY (consumer_axi_gp5_awready),
.SAXIGP5WDATA (consumer_axi_gp5_wdata),
.SAXIGP5WSTRB (consumer_axi_gp5_wstrb),
.SAXIGP5WLAST (consumer_axi_gp5_wlast),
.SAXIGP5WVALID (consumer_axi_gp5_wvalid),
.SAXIGP5WREADY (consumer_axi_gp5_wready),
.SAXIGP5BID (consumer_axi_gp5_bid),
.SAXIGP5BRESP (consumer_axi_gp5_bresp),
.SAXIGP5BVALID (consumer_axi_gp5_bvalid),
.SAXIGP5BREADY (consumer_axi_gp5_bready),
.SAXIGP5ARID (consumer_axi_gp5_arid),
.SAXIGP5ARADDR (consumer_axi_gp5_araddr),
.SAXIGP5ARLEN (consumer_axi_gp5_arlen),
.SAXIGP5ARSIZE (consumer_axi_gp5_arsize),
.SAXIGP5ARBURST (consumer_axi_gp5_arburst),
.SAXIGP5ARLOCK (consumer_axi_gp5_arlock),
.SAXIGP5ARCACHE (consumer_axi_gp5_arcache),
.SAXIGP5ARPROT (consumer_axi_gp5_arprot),
.SAXIGP5ARVALID (consumer_axi_gp5_arvalid),
.SAXIGP5ARREADY (consumer_axi_gp5_arready),
.SAXIGP5RID (consumer_axi_gp5_rid),
.SAXIGP5RDATA (consumer_axi_gp5_rdata),
.SAXIGP5RRESP (consumer_axi_gp5_rresp),
.SAXIGP5RLAST (consumer_axi_gp5_rlast),
.SAXIGP5RVALID (consumer_axi_gp5_rvalid),
.SAXIGP5RREADY (consumer_axi_gp5_rready),
.SAXIGP5AWQOS (consumer_axi_gp5_awqos),
.SAXIGP5ARQOS (consumer_axi_gp5_arqos),
.SAXIGP5RCOUNT (consumer_axi_gp5_rcount),
.SAXIGP5WCOUNT (consumer_axi_gp5_wcount),
.SAXIGP5RACOUNT (consumer_axi_gp5_racount),
.SAXIGP5WACOUNT (consumer_axi_gp5_wacount),
.SAXIGP6RCLK (clk_tps_fpl_consumer_axi_lpd_read),
.SAXIGP6WCLK (clk_tps_fpl_consumer_axi_lpd_write),
.SAXIGP6ARUSER (consumer_axi_gp6_aruser),
.SAXIGP6AWUSER (consumer_axi_gp6_awuser),
.SAXIGP6AWID (consumer_axi_gp6_awid),
.SAXIGP6AWADDR (consumer_axi_gp6_awaddr),
.SAXIGP6AWLEN (consumer_axi_gp6_awlen),
.SAXIGP6AWSIZE (consumer_axi_gp6_awsize),
.SAXIGP6AWBURST (consumer_axi_gp6_awburst),
.SAXIGP6AWLOCK (consumer_axi_gp6_awlock),
.SAXIGP6AWCACHE (consumer_axi_gp6_awcache),
.SAXIGP6AWPROT (consumer_axi_gp6_awprot),
.SAXIGP6AWVALID (consumer_axi_gp6_awvalid),
.SAXIGP6AWREADY (consumer_axi_gp6_awready),
.SAXIGP6WDATA (consumer_axi_gp6_wdata),
.SAXIGP6WSTRB (consumer_axi_gp6_wstrb),
.SAXIGP6WLAST (consumer_axi_gp6_wlast),
.SAXIGP6WVALID (consumer_axi_gp6_wvalid),
.SAXIGP6WREADY (consumer_axi_gp6_wready),
.SAXIGP6BID (consumer_axi_gp6_bid),
.SAXIGP6BRESP (consumer_axi_gp6_bresp),
.SAXIGP6BVALID (consumer_axi_gp6_bvalid),
.SAXIGP6BREADY (consumer_axi_gp6_bready),
.SAXIGP6ARID (consumer_axi_gp6_arid),
.SAXIGP6ARADDR (consumer_axi_gp6_araddr),
.SAXIGP6ARLEN (consumer_axi_gp6_arlen),
.SAXIGP6ARSIZE (consumer_axi_gp6_arsize),
.SAXIGP6ARBURST (consumer_axi_gp6_arburst),
.SAXIGP6ARLOCK (consumer_axi_gp6_arlock),
.SAXIGP6ARCACHE (consumer_axi_gp6_arcache),
.SAXIGP6ARPROT (consumer_axi_gp6_arprot),
.SAXIGP6ARVALID (consumer_axi_gp6_arvalid),
.SAXIGP6ARREADY (consumer_axi_gp6_arready),
.SAXIGP6RID (consumer_axi_gp6_rid),
.SAXIGP6RDATA (consumer_axi_gp6_rdata),
.SAXIGP6RRESP (consumer_axi_gp6_rresp),
.SAXIGP6RLAST (consumer_axi_gp6_rlast),
.SAXIGP6RVALID (consumer_axi_gp6_rvalid),
.SAXIGP6RREADY (consumer_axi_gp6_rready),
.SAXIGP6AWQOS (consumer_axi_gp6_awqos),
.SAXIGP6ARQOS (consumer_axi_gp6_arqos),
.SAXIGP6RCOUNT (consumer_axi_gp6_rcount),
.SAXIGP6WCOUNT (consumer_axi_gp6_wcount),
.SAXIGP6RACOUNT (consumer_axi_gp6_racount),
.SAXIGP6WACOUNT (consumer_axi_gp6_wacount),
.SAXIACPACLK (clk_tps_fpl_consumer_acp_fpd),
.SAXIACPAWADDR (consumer_axi_acp_awaddr),
.SAXIACPAWID (consumer_axi_acp_awid),
.SAXIACPAWLEN (consumer_axi_acp_awlen),
.SAXIACPAWSIZE (consumer_axi_acp_awsize),
.SAXIACPAWBURST (consumer_axi_acp_awburst),
.SAXIACPAWLOCK (consumer_axi_acp_awlock),
.SAXIACPAWCACHE (consumer_axi_acp_awcache),
.SAXIACPAWPROT (consumer_axi_acp_awprot),
.SAXIACPAWVALID (consumer_axi_acp_awvalid),
.SAXIACPAWREADY (consumer_axi_acp_awready),
.SAXIACPAWUSER (consumer_axi_acp_awuser),
.SAXIACPAWQOS (consumer_axi_acp_awqos),
.SAXIACPWLAST (consumer_axi_acp_wlast),
.SAXIACPWDATA (consumer_axi_acp_wdata),
.SAXIACPWSTRB (consumer_axi_acp_wstrb),
.SAXIACPWVALID (consumer_axi_acp_wvalid),
.SAXIACPWREADY (consumer_axi_acp_wready),
.SAXIACPBRESP (consumer_axi_acp_bresp),
.SAXIACPBID (consumer_axi_acp_bid),
.SAXIACPBVALID (consumer_axi_acp_bvalid),
.SAXIACPBREADY (consumer_axi_acp_bready),
.SAXIACPARADDR (consumer_axi_acp_araddr),
.SAXIACPARID (consumer_axi_acp_arid),
.SAXIACPARLEN (consumer_axi_acp_arlen),
.SAXIACPARSIZE (consumer_axi_acp_arsize),
.SAXIACPARBURST (consumer_axi_acp_arburst),
.SAXIACPARLOCK (consumer_axi_acp_arlock),
.SAXIACPARCACHE (consumer_axi_acp_arcache),
.SAXIACPARPROT (consumer_axi_acp_arprot),
.SAXIACPARVALID (consumer_axi_acp_arvalid),
.SAXIACPARREADY (consumer_axi_acp_arready),
.SAXIACPARUSER (consumer_axi_acp_aruser),
.SAXIACPARQOS (consumer_axi_acp_arqos),
.SAXIACPRID (consumer_axi_acp_rid),
.SAXIACPRLAST (consumer_axi_acp_rlast),
.SAXIACPRDATA (consumer_axi_acp_rdata),
.SAXIACPRRESP (consumer_axi_acp_rresp),
.SAXIACPRVALID (consumer_axi_acp_rvalid),
.SAXIACPRREADY (consumer_axi_acp_rready),
.PLACECLK (consumer_axi_ace_fpd_aclk),
.SACEFPDAWVALID (consumer_axi_ace_fpd_awvalid),
.SACEFPDAWREADY (consumer_axi_ace_fpd_awready),
.SACEFPDAWID (consumer_axi_ace_fpd_awid),
.SACEFPDAWADDR (consumer_axi_ace_fpd_awaddr),
.SACEFPDAWREGION (consumer_axi_ace_fpd_awregion),
.SACEFPDAWLEN (consumer_axi_ace_fpd_awlen),
.SACEFPDAWSIZE (consumer_axi_ace_fpd_awsize),
.SACEFPDAWBURST (consumer_axi_ace_fpd_awburst),
.SACEFPDAWLOCK (consumer_axi_ace_fpd_awlock),
.SACEFPDAWCACHE (consumer_axi_ace_fpd_awcache),
.SACEFPDAWPROT (consumer_axi_ace_fpd_awprot),
.SACEFPDAWDOMAIN (consumer_axi_ace_fpd_awdomain),
.SACEFPDAWSNOOP (consumer_axi_ace_fpd_awsnoop),
.SACEFPDAWBAR (consumer_axi_ace_fpd_awbar),
.SACEFPDAWQOS (consumer_axi_ace_fpd_awqos),
.SACEFPDAWUSER (consumer_axi_ace_fpd_awuser),
.SACEFPDWVALID (consumer_axi_ace_fpd_wvalid),
.SACEFPDWREADY (consumer_axi_ace_fpd_wready),
.SACEFPDWDATA (consumer_axi_ace_fpd_wdata),
.SACEFPDWSTRB (consumer_axi_ace_fpd_wstrb),
.SACEFPDWLAST (consumer_axi_ace_fpd_wlast),
.SACEFPDWUSER (consumer_axi_ace_fpd_wuser),
.SACEFPDBVALID (consumer_axi_ace_fpd_bvalid),
.SACEFPDBREADY (consumer_axi_ace_fpd_bready),
.SACEFPDBID (consumer_axi_ace_fpd_bid),
.SACEFPDBRESP (consumer_axi_ace_fpd_bresp),
.SACEFPDBUSER (consumer_axi_ace_fpd_buser),
.SACEFPDARVALID (consumer_axi_ace_fpd_arvalid),
.SACEFPDARREADY (consumer_axi_ace_fpd_arready),
.SACEFPDARID (consumer_axi_ace_fpd_arid),
.SACEFPDARADDR (consumer_axi_ace_fpd_araddr),
.SACEFPDARREGION (consumer_axi_ace_fpd_arregion),
.SACEFPDARLEN (consumer_axi_ace_fpd_arlen),
.SACEFPDARSIZE (consumer_axi_ace_fpd_arsize),
.SACEFPDARBURST (consumer_axi_ace_fpd_arburst),
.SACEFPDARLOCK (consumer_axi_ace_fpd_arlock),
.SACEFPDARCACHE (consumer_axi_ace_fpd_arcache),
.SACEFPDARPROT (consumer_axi_ace_fpd_arprot),
.SACEFPDARDOMAIN (consumer_axi_ace_fpd_ardomain),
.SACEFPDARSNOOP (consumer_axi_ace_fpd_arsnoop),
.SACEFPDARBAR (consumer_axi_ace_fpd_arbar),
.SACEFPDARQOS (consumer_axi_ace_fpd_arqos),
.SACEFPDARUSER (consumer_axi_ace_fpd_aruser),
.SACEFPDRVALID (consumer_axi_ace_fpd_rvalid),
.SACEFPDRREADY (consumer_axi_ace_fpd_rready),
.SACEFPDRID (consumer_axi_ace_fpd_rid),
.SACEFPDRDATA (consumer_axi_ace_fpd_rdata),
.SACEFPDRRESP (consumer_axi_ace_fpd_rresp),
.SACEFPDRLAST (consumer_axi_ace_fpd_rlast),
.SACEFPDRUSER (consumer_axi_ace_fpd_ruser),
.SACEFPDACVALID (consumer_axi_ace_fpd_acvalid),
.SACEFPDACREADY (consumer_axi_ace_fpd_acready),
.SACEFPDACADDR (consumer_axi_ace_fpd_acaddr),
.SACEFPDACSNOOP (consumer_axi_ace_fpd_acsnoop),
.SACEFPDACPROT (consumer_axi_ace_fpd_acprot),
.SACEFPDCRVALID (consumer_axi_ace_fpd_crvalid),
.SACEFPDCRREADY (consumer_axi_ace_fpd_crready),
.SACEFPDCRRESP (consumer_axi_ace_fpd_crresp),
.SACEFPDCDVALID (consumer_axi_ace_fpd_cdvalid),
.SACEFPDCDREADY (consumer_axi_ace_fpd_cdready),
.SACEFPDCDDATA (consumer_axi_ace_fpd_cddata),
.SACEFPDCDLAST (consumer_axi_ace_fpd_cdlast),
.SACEFPDWACK (consumer_axi_ace_fpd_wack),
.SACEFPDRACK (consumer_axi_ace_fpd_rack),
.EMIOCAN0PHYTX (emio_can0_phy_tx),
.EMIOCAN0PHYRX (emio_can0_phy_rx),
.EMIOCAN1PHYTX (emio_can1_phy_tx),
.EMIOCAN1PHYRX (emio_can1_phy_rx),
.EMIOENET0GMIIRXCLK (clk_tps_fpl_emio_enet0_gmii_rx),
.EMIOENET0SPEEDMODE (emio_enet0_speed_mode),
.EMIOENET0GMIICRS (emio_enet0_gmii_crs),
.EMIOENET0GMIICOL (emio_enet0_gmii_col),
.EMIOENET0GMIIRXD (emio_enet0_gmii_rxd),
.EMIOENET0GMIIRXER (emio_enet0_gmii_rx_er),
.EMIOENET0GMIIRXDV (emio_enet0_gmii_rx_dv),
.EMIOENET0GMIITXCLK (clk_tps_fpl_emio_enet0_gmii_tx),
.EMIOENET0GMIITXD (emio_enet0_gmii_txd),
.EMIOENET0GMIITXEN (emio_enet0_gmii_tx_en),
.EMIOENET0GMIITXER (emio_enet0_gmii_tx_er),
.EMIOENET0MDIOMDC (emio_enet0_mdio_mdc),
.EMIOENET0MDIOI (emio_enet0_mdio_i),
.EMIOENET0MDIOO (emio_enet0_mdio_o),
.EMIOENET0MDIOTN (emio_enet0_mdio_t_n),
.EMIOENET1GMIIRXCLK (clk_tps_fpl_emio_enet1_gmii_rx),
.EMIOENET1SPEEDMODE (emio_enet1_speed_mode),
.EMIOENET1GMIICRS (emio_enet1_gmii_crs),
.EMIOENET1GMIICOL (emio_enet1_gmii_col),
.EMIOENET1GMIIRXD (emio_enet1_gmii_rxd),
.EMIOENET1GMIIRXER (emio_enet1_gmii_rx_er),
.EMIOENET1GMIIRXDV (emio_enet1_gmii_rx_dv),
.EMIOENET1GMIITXCLK (clk_tps_fpl_emio_enet1_gmii_tx),
.EMIOENET1GMIITXD (emio_enet1_gmii_txd),
.EMIOENET1GMIITXEN (emio_enet1_gmii_tx_en),
.EMIOENET1GMIITXER (emio_enet1_gmii_tx_er),
.EMIOENET1MDIOMDC (emio_enet1_mdio_mdc),
.EMIOENET1MDIOI (emio_enet1_mdio_i),
.EMIOENET1MDIOO (emio_enet1_mdio_o),
.EMIOENET1MDIOTN (emio_enet1_mdio_t_n),
.EMIOENET2GMIIRXCLK (clk_tps_fpl_emio_enet2_gmii_rx),
.EMIOENET2SPEEDMODE (emio_enet2_speed_mode),
.EMIOENET2GMIICRS (emio_enet2_gmii_crs),
.EMIOENET2GMIICOL (emio_enet2_gmii_col),
.EMIOENET2GMIIRXD (emio_enet2_gmii_rxd),
.EMIOENET2GMIIRXER (emio_enet2_gmii_rx_er),
.EMIOENET2GMIIRXDV (emio_enet2_gmii_rx_dv),
.EMIOENET2GMIITXCLK (clk_tps_fpl_emio_enet2_gmii_tx),
.EMIOENET2GMIITXD (emio_enet2_gmii_txd),
.EMIOENET2GMIITXEN (emio_enet2_gmii_tx_en),
.EMIOENET2GMIITXER (emio_enet2_gmii_tx_er),
.EMIOENET2MDIOMDC (emio_enet2_mdio_mdc),
.EMIOENET2MDIOI (emio_enet2_mdio_i),
.EMIOENET2MDIOO (emio_enet2_mdio_o),
.EMIOENET2MDIOTN (emio_enet2_mdio_t_n),
.EMIOENET3GMIIRXCLK (clk_tps_fpl_emio_enet3_gmii_rx),
.EMIOENET3SPEEDMODE (emio_enet3_speed_mode),
.EMIOENET3GMIICRS (emio_enet3_gmii_crs),
.EMIOENET3GMIICOL (emio_enet3_gmii_col),
.EMIOENET3GMIIRXD (emio_enet3_gmii_rxd),
.EMIOENET3GMIIRXER (emio_enet3_gmii_rx_er),
.EMIOENET3GMIIRXDV (emio_enet3_gmii_rx_dv),
.EMIOENET3GMIITXCLK (clk_tps_fpl_emio_enet3_gmii_tx),
.EMIOENET3GMIITXD (emio_enet3_gmii_txd),
.EMIOENET3GMIITXEN (emio_enet3_gmii_tx_en),
.EMIOENET3GMIITXER (emio_enet3_gmii_tx_er),
.EMIOENET3MDIOMDC (emio_enet3_mdio_mdc),
.EMIOENET3MDIOI (emio_enet3_mdio_i),
.EMIOENET3MDIOO (emio_enet3_mdio_o),
.EMIOENET3MDIOTN (emio_enet3_mdio_t_n),
.EMIOENET0TXRDATARDY (emio_enet0_tx_r_data_rdy),
.EMIOENET0TXRRD (emio_enet0_tx_r_rd),
.EMIOENET0TXRVALID (emio_enet0_tx_r_valid),
.EMIOENET0TXRDATA (emio_enet0_tx_r_data),
.EMIOENET0TXRSOP (emio_enet0_tx_r_sop),
.EMIOENET0TXREOP (emio_enet0_tx_r_eop),
.EMIOENET0TXRERR (emio_enet0_tx_r_err),
.EMIOENET0TXRUNDERFLOW (emio_enet0_tx_r_underflow),
.EMIOENET0TXRFLUSHED (emio_enet0_tx_r_flushed),
.EMIOENET0TXRCONTROL (emio_enet0_tx_r_control),
.EMIOENET0DMATXENDTOG (emio_enet0_dma_tx_end_tog),
.EMIOENET0DMATXSTATUSTOG (emio_enet0_dma_tx_status_tog),
.EMIOENET0TXRSTATUS (emio_enet0_tx_r_status),
.EMIOENET0RXWWR (emio_enet0_rx_w_wr),
.EMIOENET0RXWDATA (emio_enet0_rx_w_data),
.EMIOENET0RXWSOP (emio_enet0_rx_w_sop),
.EMIOENET0RXWEOP (emio_enet0_rx_w_eop),
.EMIOENET0RXWSTATUS (emio_enet0_rx_w_status),
.EMIOENET0RXWERR (emio_enet0_rx_w_err),
.EMIOENET0RXWOVERFLOW (emio_enet0_rx_w_overflow),
.FMIOGEM0SIGNALDETECT (emio_enet0_signal_detect),
.EMIOENET0RXWFLUSH (emio_enet0_rx_w_flush),
.EMIOGEM0TXRFIXEDLAT (emio_enet0_tx_r_fixed_lat),
.FMIOGEM0FIFOTXCLKFROMPL (clk_tps_fpl_fmio_gem0_fifo_tx),
.FMIOGEM0FIFORXCLKFROMPL (clk_tps_fpl_fmio_gem0_fifo_rx),
.FMIOGEM0FIFOTXCLKTOPLBUFG (clk_fps_tpl_fmio_gem0_fifo_tx),
.FMIOGEM0FIFORXCLKTOPLBUFG (clk_fps_tpl_fmio_gem0_fifo_rx),
.EMIOENET1TXRDATARDY (emio_enet1_tx_r_data_rdy),
.EMIOENET1TXRRD (emio_enet1_tx_r_rd),
.EMIOENET1TXRVALID (emio_enet1_tx_r_valid),
.EMIOENET1TXRDATA (emio_enet1_tx_r_data),
.EMIOENET1TXRSOP (emio_enet1_tx_r_sop),
.EMIOENET1TXREOP (emio_enet1_tx_r_eop),
.EMIOENET1TXRERR (emio_enet1_tx_r_err),
.EMIOENET1TXRUNDERFLOW (emio_enet1_tx_r_underflow),
.EMIOENET1TXRFLUSHED (emio_enet1_tx_r_flushed),
.EMIOENET1TXRCONTROL (emio_enet1_tx_r_control),
.EMIOENET1DMATXENDTOG (emio_enet1_dma_tx_end_tog),
.EMIOENET1DMATXSTATUSTOG (emio_enet1_dma_tx_status_tog),
.EMIOENET1TXRSTATUS (emio_enet1_tx_r_status),
.EMIOENET1RXWWR (emio_enet1_rx_w_wr),
.EMIOENET1RXWDATA (emio_enet1_rx_w_data),
.EMIOENET1RXWSOP (emio_enet1_rx_w_sop),
.EMIOENET1RXWEOP (emio_enet1_rx_w_eop),
.EMIOENET1RXWSTATUS (emio_enet1_rx_w_status),
.EMIOENET1RXWERR (emio_enet1_rx_w_err),
.EMIOENET1RXWOVERFLOW (emio_enet1_rx_w_overflow),
.FMIOGEM1SIGNALDETECT (emio_enet1_signal_detect),
.EMIOENET1RXWFLUSH (emio_enet1_rx_w_flush),
.EMIOGEM1TXRFIXEDLAT (emio_enet1_tx_r_fixed_lat),
.FMIOGEM1FIFOTXCLKFROMPL (clk_tps_fpl_fmio_gem1_fifo_tx),
.FMIOGEM1FIFORXCLKFROMPL (clk_tps_fpl_fmio_gem1_fifo_rx),
.FMIOGEM1FIFOTXCLKTOPLBUFG (clk_fps_tpl_fmio_gem1_fifo_tx),
.FMIOGEM1FIFORXCLKTOPLBUFG (clk_fps_tpl_fmio_gem1_fifo_rx),
.EMIOENET2TXRDATARDY (emio_enet2_tx_r_data_rdy),
.EMIOENET2TXRRD (emio_enet2_tx_r_rd),
.EMIOENET2TXRVALID (emio_enet2_tx_r_valid),
.EMIOENET2TXRDATA (emio_enet2_tx_r_data),
.EMIOENET2TXRSOP (emio_enet2_tx_r_sop),
.EMIOENET2TXREOP (emio_enet2_tx_r_eop),
.EMIOENET2TXRERR (emio_enet2_tx_r_err),
.EMIOENET2TXRUNDERFLOW (emio_enet2_tx_r_underflow),
.EMIOENET2TXRFLUSHED (emio_enet2_tx_r_flushed),
.EMIOENET2TXRCONTROL (emio_enet2_tx_r_control),
.EMIOENET2DMATXENDTOG (emio_enet2_dma_tx_end_tog),
.EMIOENET2DMATXSTATUSTOG (emio_enet2_dma_tx_status_tog),
.EMIOENET2TXRSTATUS (emio_enet2_tx_r_status),
.EMIOENET2RXWWR (emio_enet2_rx_w_wr),
.EMIOENET2RXWDATA (emio_enet2_rx_w_data),
.EMIOENET2RXWSOP (emio_enet2_rx_w_sop),
.EMIOENET2RXWEOP (emio_enet2_rx_w_eop),
.EMIOENET2RXWSTATUS (emio_enet2_rx_w_status),
.EMIOENET2RXWERR (emio_enet2_rx_w_err),
.EMIOENET2RXWOVERFLOW (emio_enet2_rx_w_overflow),
.FMIOGEM2SIGNALDETECT (emio_enet2_signal_detect),
.EMIOENET2RXWFLUSH (emio_enet2_rx_w_flush),
.EMIOGEM2TXRFIXEDLAT (emio_enet2_tx_r_fixed_lat),
.FMIOGEM2FIFOTXCLKFROMPL (clk_tps_fpl_fmio_gem2_fifo_tx),
.FMIOGEM2FIFORXCLKFROMPL (clk_tps_fpl_fmio_gem2_fifo_rx),
.FMIOGEM2FIFOTXCLKTOPLBUFG (clk_fps_tpl_fmio_gem2_fifo_tx),
.FMIOGEM2FIFORXCLKTOPLBUFG (clk_fps_tpl_fmio_gem2_fifo_rx),
.EMIOENET3TXRDATARDY (emio_enet3_tx_r_data_rdy),
.EMIOENET3TXRRD (emio_enet3_tx_r_rd),
.EMIOENET3TXRVALID (emio_enet3_tx_r_valid),
.EMIOENET3TXRDATA (emio_enet3_tx_r_data),
.EMIOENET3TXRSOP (emio_enet3_tx_r_sop),
.EMIOENET3TXREOP (emio_enet3_tx_r_eop),
.EMIOENET3TXRERR (emio_enet3_tx_r_err),
.EMIOENET3TXRUNDERFLOW (emio_enet3_tx_r_underflow),
.EMIOENET3TXRFLUSHED (emio_enet3_tx_r_flushed),
.EMIOENET3TXRCONTROL (emio_enet3_tx_r_control),
.EMIOENET3DMATXENDTOG (emio_enet3_dma_tx_end_tog),
.EMIOENET3DMATXSTATUSTOG (emio_enet3_dma_tx_status_tog),
.EMIOENET3TXRSTATUS (emio_enet3_tx_r_status),
.EMIOENET3RXWWR (emio_enet3_rx_w_wr),
.EMIOENET3RXWDATA (emio_enet3_rx_w_data),
.EMIOENET3RXWSOP (emio_enet3_rx_w_sop),
.EMIOENET3RXWEOP (emio_enet3_rx_w_eop),
.EMIOENET3RXWSTATUS (emio_enet3_rx_w_status),
.EMIOENET3RXWERR (emio_enet3_rx_w_err),
.EMIOENET3RXWOVERFLOW (emio_enet3_rx_w_overflow),
.FMIOGEM3SIGNALDETECT (emio_enet3_signal_detect),
.EMIOENET3RXWFLUSH (emio_enet3_rx_w_flush),
.EMIOGEM3TXRFIXEDLAT (emio_enet3_tx_r_fixed_lat),
.FMIOGEM3FIFOTXCLKFROMPL (clk_tps_fpl_fmio_gem3_fifo_tx),
.FMIOGEM3FIFORXCLKFROMPL (clk_tps_fpl_fmio_gem3_fifo_rx),
.FMIOGEM3FIFOTXCLKTOPLBUFG (clk_fps_tpl_fmio_gem3_fifo_tx),
.FMIOGEM3FIFORXCLKTOPLBUFG (clk_fps_tpl_fmio_gem3_fifo_rx),
.EMIOGEM0TXSOF (emio_enet0_tx_sof),
.EMIOGEM0SYNCFRAMETX (emio_enet0_sync_frame_tx),
.EMIOGEM0DELAYREQTX (emio_enet0_delay_req_tx),
.EMIOGEM0PDELAYREQTX (emio_enet0_pdelay_req_tx),
.EMIOGEM0PDELAYRESPTX (emio_enet0_pdelay_resp_tx),
.EMIOGEM0RXSOF (emio_enet0_rx_sof),
.EMIOGEM0SYNCFRAMERX (emio_enet0_sync_frame_rx),
.EMIOGEM0DELAYREQRX (emio_enet0_delay_req_rx),
.EMIOGEM0PDELAYREQRX (emio_enet0_pdelay_req_rx),
.EMIOGEM0PDELAYRESPRX (emio_enet0_pdelay_resp_rx),
.EMIOGEM0TSUINCCTRL (emio_enet0_tsu_inc_ctrl),
.EMIOGEM0TSUTIMERCMPVAL (emio_enet0_tsu_timer_cmp_val),
.EMIOGEM1TXSOF (emio_enet1_tx_sof),
.EMIOGEM1SYNCFRAMETX (emio_enet1_sync_frame_tx),
.EMIOGEM1DELAYREQTX (emio_enet1_delay_req_tx),
.EMIOGEM1PDELAYREQTX (emio_enet1_pdelay_req_tx),
.EMIOGEM1PDELAYRESPTX (emio_enet1_pdelay_resp_tx),
.EMIOGEM1RXSOF (emio_enet1_rx_sof),
.EMIOGEM1SYNCFRAMERX (emio_enet1_sync_frame_rx),
.EMIOGEM1DELAYREQRX (emio_enet1_delay_req_rx),
.EMIOGEM1PDELAYREQRX (emio_enet1_pdelay_req_rx),
.EMIOGEM1PDELAYRESPRX (emio_enet1_pdelay_resp_rx),
.EMIOGEM1TSUINCCTRL (emio_enet1_tsu_inc_ctrl),
.EMIOGEM1TSUTIMERCMPVAL (emio_enet1_tsu_timer_cmp_val),
.EMIOGEM2TXSOF (emio_enet2_tx_sof),
.EMIOGEM2SYNCFRAMETX (emio_enet2_sync_frame_tx),
.EMIOGEM2DELAYREQTX (emio_enet2_delay_req_tx),
.EMIOGEM2PDELAYREQTX (emio_enet2_pdelay_req_tx),
.EMIOGEM2PDELAYRESPTX (emio_enet2_pdelay_resp_tx),
.EMIOGEM2RXSOF (emio_enet2_rx_sof),
.EMIOGEM2SYNCFRAMERX (emio_enet2_sync_frame_rx),
.EMIOGEM2DELAYREQRX (emio_enet2_delay_req_rx),
.EMIOGEM2PDELAYREQRX (emio_enet2_pdelay_req_rx),
.EMIOGEM2PDELAYRESPRX (emio_enet2_pdelay_resp_rx),
.EMIOGEM2TSUINCCTRL (emio_enet2_tsu_inc_ctrl),
.EMIOGEM2TSUTIMERCMPVAL (emio_enet2_tsu_timer_cmp_val),
.EMIOGEM3TXSOF (emio_enet3_tx_sof),
.EMIOGEM3SYNCFRAMETX (emio_enet3_sync_frame_tx),
.EMIOGEM3DELAYREQTX (emio_enet3_delay_req_tx),
.EMIOGEM3PDELAYREQTX (emio_enet3_pdelay_req_tx),
.EMIOGEM3PDELAYRESPTX (emio_enet3_pdelay_resp_tx),
.EMIOGEM3RXSOF (emio_enet3_rx_sof),
.EMIOGEM3SYNCFRAMERX (emio_enet3_sync_frame_rx),
.EMIOGEM3DELAYREQRX (emio_enet3_delay_req_rx),
.EMIOGEM3PDELAYREQRX (emio_enet3_pdelay_req_rx),
.EMIOGEM3PDELAYRESPRX (emio_enet3_pdelay_resp_rx),
.EMIOGEM3TSUINCCTRL (emio_enet3_tsu_inc_ctrl),
.EMIOGEM3TSUTIMERCMPVAL (emio_enet3_tsu_timer_cmp_val),
.FMIOGEMTSUCLKFROMPL (clk_tps_fpl_fmio_gem_tsu),
.FMIOGEMTSUCLKTOPLBUFG (clk_fps_tpl_gem_tsu_clk),
.EMIOENETTSUCLK (clk_tps_fpl_emio_enet_tsu),
.EMIOENET0GEMTSUTIMERCNT (emio_enet0_enet_tsu_timer_cnt),
.EMIOENET0EXTINTIN (emio_enet0_ext_int_in),
.EMIOENET1EXTINTIN (emio_enet1_ext_int_in),
.EMIOENET2EXTINTIN (emio_enet2_ext_int_in),
.EMIOENET3EXTINTIN (emio_enet3_ext_int_in),
.EMIOENET0DMABUSWIDTH (emio_enet0_dma_bus_width),
.EMIOENET1DMABUSWIDTH (emio_enet1_dma_bus_width),
.EMIOENET2DMABUSWIDTH (emio_enet2_dma_bus_width),
.EMIOENET3DMABUSWIDTH (emio_enet3_dma_bus_width),
.EMIOGPIOI (emio_gpio_i),
.EMIOGPIOO (emio_gpio_o),
.EMIOGPIOTN (emio_gpio_t_n),
.EMIOI2C0SCLI (emio_i2c0_scl_i),
.EMIOI2C0SCLO (emio_i2c0_scl_o),
.EMIOI2C0SCLTN (emio_i2c0_scl_tri),
.EMIOI2C0SDAI (emio_i2c0_sda_i),
.EMIOI2C0SDAO (emio_i2c0_sda_o),
.EMIOI2C0SDATN (emio_i2c0_sda_t_n),
.EMIOI2C1SCLI (emio_i2c1_scl_i),
.EMIOI2C1SCLO (emio_i2c1_scl_o),
.EMIOI2C1SCLTN (emio_i2c1_scl_tri),
.EMIOI2C1SDAI (emio_i2c1_sda_i),
.EMIOI2C1SDAO (emio_i2c1_sda_o),
.EMIOI2C1SDATN (emio_i2c1_sda_t_n),
.EMIOUART0TX (emio_uart0_txd),
.EMIOUART0RX (emio_uart0_rxd),
.EMIOUART0CTSN (emio_uart0_ctsn),
.EMIOUART0RTSN (emio_uart0_rtsn),
.EMIOUART0DSRN (emio_uart0_dsrn),
.EMIOUART0DCDN (emio_uart0_dcdn),
.EMIOUART0RIN (emio_uart0_rin),
.EMIOUART0DTRN (emio_uart0_dtrn),
.EMIOUART1TX (emio_uart1_txd),
.EMIOUART1RX (emio_uart1_rxd),
.EMIOUART1CTSN (emio_uart1_ctsn),
.EMIOUART1RTSN (emio_uart1_rtsn),
.EMIOUART1DSRN (emio_uart1_dsrn),
.EMIOUART1DCDN (emio_uart1_dcdn),
.EMIOUART1RIN (emio_uart1_rin),
.EMIOUART1DTRN (emio_uart1_dtrn),
.EMIOSDIO0CLKOUT (clk_fps_tpl_emio_sdio0),
.EMIOSDIO0FBCLKIN (clk_tps_fpl_emio_sdio0),
.EMIOSDIO0CMDOUT (emio_sdio0_cmdout),
.EMIOSDIO0CMDIN (emio_sdio0_cmdin),
.EMIOSDIO0CMDENA (emio_sdio0_cmdena_n),
.EMIOSDIO0DATAIN (emio_sdio0_datain),
.EMIOSDIO0DATAOUT (emio_sdio0_dataout),
.EMIOSDIO0DATAENA (emio_sdio0_dataena_n),
.EMIOSDIO0CDN (emio_sdio0_cd_n),
.EMIOSDIO0WP (emio_sdio0_wp),
.EMIOSDIO0LEDCONTROL (emio_sdio0_ledcontrol),
.EMIOSDIO0BUSPOWER (emio_sdio0_buspower),
.EMIOSDIO0BUSVOLT (emio_sdio0_bus_volt),
.EMIOSDIO1CLKOUT (clk_fps_tpl_emio_sdio1),
.EMIOSDIO1FBCLKIN (clk_tps_fpl_emio_sdio1),
.EMIOSDIO1CMDOUT (emio_sdio1_cmdout),
.EMIOSDIO1CMDIN (emio_sdio1_cmdin),
.EMIOSDIO1CMDENA (emio_sdio1_cmdena_n),
.EMIOSDIO1DATAIN (emio_sdio1_datain),
.EMIOSDIO1DATAOUT (emio_sdio1_dataout),
.EMIOSDIO1DATAENA (emio_sdio1_dataena_n),
.EMIOSDIO1CDN (emio_sdio1_cd_n),
.EMIOSDIO1WP (emio_sdio1_wp),
.EMIOSDIO1LEDCONTROL (emio_sdio1_ledcontrol),
.EMIOSDIO1BUSPOWER (emio_sdio1_buspower),
.EMIOSDIO1BUSVOLT (emio_sdio1_bus_volt),
.EMIOSPI0SCLKI (emio_spi0_sclk_i),
.EMIOSPI0SCLKO (emio_spi0_sclk_o),
.EMIOSPI0SCLKTN (emio_spi0_sclk_t_n),
.EMIOSPI0MI (emio_spi0_m_i),
.EMIOSPI0MO (emio_spi0_m_o),
.EMIOSPI0MOTN (emio_spi0_mo_t_n),
.EMIOSPI0SI (emio_spi0_s_i),
.EMIOSPI0SO (emio_spi0_s_o),
.EMIOSPI0STN (emio_spi0_so_t_n),
.EMIOSPI0SSIN (emio_spi0_ss_i_n),
.EMIOSPI0SSON ({emio_spi0_ss2_o_n,emio_spi0_ss1_o_n,emio_spi0_ss_o_n}),
.EMIOSPI0SSNTN (emio_spi0_ss_n_t_n),
.EMIOSPI1SCLKI (emio_spi1_sclk_i),
.EMIOSPI1SCLKO (emio_spi1_sclk_o),
.EMIOSPI1SCLKTN (emio_spi1_sclk_t_n),
.EMIOSPI1MI (emio_spi1_m_i),
.EMIOSPI1MO (emio_spi1_m_o),
.EMIOSPI1MOTN (emio_spi1_mo_t_n),
.EMIOSPI1SI (emio_spi1_s_i),
.EMIOSPI1SO (emio_spi1_s_o),
.EMIOSPI1STN (emio_spi1_so_tri),
.EMIOSPI1SSIN (emio_spi1_ss_i_n),
.EMIOSPI1SSON ({emio_spi1_ss2_o_n,emio_spi1_ss1_o_n,emio_spi1_ss_o_n}),
.EMIOSPI1SSNTN (emio_spi1_ss_n_t_n),
.PLPSTRACECLK (clk_tps_fpl_trace),
.PSPLTRACECTL (ps_pl_tracectl),
.PSPLTRACEDATA (ps_pl_tracedata),
.EMIOTTC0WAVEO (emio_ttc0_wave_o),
.EMIOTTC0CLKI (clk_tps_fpl_emio_ttc0),
.EMIOTTC1WAVEO (emio_ttc1_wave_o),
.EMIOTTC1CLKI (clk_tps_fpl_emio_ttc1),
.EMIOTTC2WAVEO (emio_ttc2_wave_o),
.EMIOTTC2CLKI (clk_tps_fpl_emio_ttc2),
.EMIOTTC3WAVEO (emio_ttc3_wave_o),
.EMIOTTC3CLKI (clk_tps_fpl_emio_ttc3),
.EMIOWDT0CLKI (clk_tps_fpl_emio_wdt0),
.EMIOWDT0RSTO (emio_wdt0_rst_o),
.EMIOWDT1CLKI (clk_tps_fpl_emio_wdt1),
.EMIOWDT1RSTO (emio_wdt1_rst_o),
.EMIOHUBPORTOVERCRNTUSB30 (emio_hub_port_overcrnt_usb3_0),
.EMIOHUBPORTOVERCRNTUSB31 (emio_hub_port_overcrnt_usb3_1),
.EMIOHUBPORTOVERCRNTUSB20 (emio_hub_port_overcrnt_usb2_0),
.EMIOHUBPORTOVERCRNTUSB21 (emio_hub_port_overcrnt_usb2_1),
.EMIOU2DSPORTVBUSCTRLUSB30 (emio_u2dsport_vbus_ctrl_usb3_0),
.EMIOU2DSPORTVBUSCTRLUSB31 (emio_u2dsport_vbus_ctrl_usb3_1),
.EMIOU3DSPORTVBUSCTRLUSB30 (emio_u3dsport_vbus_ctrl_usb3_0),
.EMIOU3DSPORTVBUSCTRLUSB31 (emio_u3dsport_vbus_ctrl_usb3_1),
.ADMAFCICLK (clk_tps_fpl_adma_fci),
.PL2ADMACVLD (pl2adma_cvld),
.PL2ADMATACK (pl2adma_tack),
.ADMA2PLCACK (adma2pl_cack),
.ADMA2PLTVLD (adma2pl_tvld),
.GDMAFCICLK (clk_tps_fpl_gdma_perif),
.PL2GDMACVLD (perif_gdma_cvld),
.PL2GDMATACK (perif_gdma_tack),
.GDMA2PLCACK (gdma_perif_cack),
.GDMA2PLTVLD (gdma_perif_tvld),
.PLFPGASTOP (pl_clock_stop),
.PLLAUXREFCLKLPD (clk_tps_fpl_pll_aux_lpd),
.PLLAUXREFCLKFPD (clk_tps_fpl_pll_aux_fpd),
.DPSAXISAUDIOTDATA (consumer_axi_stream_dp_audio_tdata),
.DPSAXISAUDIOTID (consumer_axi_stream_dp_audio_tid),
.DPSAXISAUDIOTVALID (consumer_axi_stream_dp_audio_tvalid),
.DPSAXISAUDIOTREADY (consumer_axi_stream_dp_audio_tready),
.DPMAXISMIXEDAUDIOTDATA (supplier_axi_stream_dp_mixed_audio_tdata),
.DPMAXISMIXEDAUDIOTID (supplier_axi_stream_dp_mixed_audio_tid),
.DPMAXISMIXEDAUDIOTVALID (supplier_axi_stream_dp_mixed_audio_tvalid),
.DPMAXISMIXEDAUDIOTREADY (supplier_axi_stream_dp_mixed_audio_tready),
.DPSAXISAUDIOCLK (clk_tps_fpl_dp_s_axis_audio),
.DPLIVEVIDEOINVSYNC (dp_live_video_in_vsync),
.DPLIVEVIDEOINHSYNC (dp_live_video_in_hsync),
.DPLIVEVIDEOINDE (dp_live_video_in_de),
.DPLIVEVIDEOINPIXEL1 (dp_live_video_in_pixel1),
.DPVIDEOINCLK (clk_tps_fpl_dp_video_in),
.DPVIDEOOUTHSYNC (dp_video_out_hsync),
.DPVIDEOOUTVSYNC (dp_video_out_vsync),
.DPVIDEOOUTPIXEL1 (dp_video_out_pixel1),
.DPAUXDATAIN (dp_aux_data_in),
.DPAUXDATAOUT (dp_aux_data_out),
.DPAUXDATAOEN (dp_aux_data_oe_n),
.DPLIVEGFXALPHAIN (dp_live_gfx_alpha_in),
.DPLIVEGFXPIXEL1IN (dp_live_gfx_pixel1_in),
.DPHOTPLUGDETECT (dp_hot_plug_detect),
.DPEXTERNALCUSTOMEVENT1 (dp_external_custom_event1),
.DPEXTERNALCUSTOMEVENT2 (dp_external_custom_event2),
.DPEXTERNALVSYNCEVENT (dp_external_vsync_event),
.DPLIVEVIDEODEOUT (dp_live_video_de_out),
.PLPSEVENTI (pl_ps_eventi),
.PSPLEVENTO (ps_pl_evento),
.PSPLSTANDBYWFE (ps_pl_standbywfe),
.PSPLSTANDBYWFI (ps_pl_standbywfi),
.PLPSAPUGICIRQ (pl_ps_apugic_irq),
.PLPSAPUGICFIQ (pl_ps_apugic_fiq),
.RPUEVENTI0 (rpu_eventi0),
.RPUEVENTI1 (rpu_eventi1),
.RPUEVENTO0 (rpu_evento0),
.RPUEVENTO1 (rpu_evento1),
.NFIQ0LPDRPU (nfiq0_lpd_rpu),
.NFIQ1LPDRPU (nfiq1_lpd_rpu),
.NIRQ0LPDRPU (nirq0_lpd_rpu),
.NIRQ1LPDRPU (nirq1_lpd_rpu),
.STMEVENT (stm_event),
.PLPSTRIGACK (pl_ps_trigack),
.PLPSTRIGGER (pl_ps_trigger),
.PSPLTRIGACK (ps_pl_trigack),
.PSPLTRIGGER (ps_pl_trigger),
.FTMGPO (ftm_gpo),
.FTMGPI (ftm_gpi),
.PLPSIRQ0 (pl_ps_irq0),
.PLPSIRQ1 (pl_ps_irq1),
.PSPLIRQLPD ({irq_lpd_dev_null[18:8],
							fps_tpl_irq_xmpu_lpd, 
							fps_tpl_irq_efuse, 
							fps_tpl_irq_csu_dma, 
							fps_tpl_irq_csu, 
							fps_tpl_irq_adma_chan, 
							fps_tpl_irq_usb3_0_pmu_wakeup, 
							fps_tpl_irq_usb3_1_otg, 
							fps_tpl_irq_usb3_1_endpoint, 
							fps_tpl_irq_usb3_0_otg, 
							fps_tpl_irq_usb3_0_endpoint, 
							fps_tpl_irq_enet3_wake, 
							fps_tpl_irq_enet3, 
							fps_tpl_irq_enet2_wake, 
							fps_tpl_irq_enet2, 
							fps_tpl_irq_enet1_wake, 
							fps_tpl_irq_enet1, 
							fps_tpl_irq_enet0_wake, 
							fps_tpl_irq_enet0, 
							fps_tpl_irq_ams, 
							fps_tpl_irq_aib_axi, 
							fps_tpl_irq_atb_err_lpd, 
							fps_tpl_irq_csu_pmu_wdt, 
							fps_tpl_irq_lp_wdt, 
							fps_tpl_irq_sdio1_wake, 
							fps_tpl_irq_sdio0_wake, 
							fps_tpl_irq_sdio1, 
							fps_tpl_irq_sdio0, 
							fps_tpl_irq_ttc3_2, 
							fps_tpl_irq_ttc3_1, 
							fps_tpl_irq_ttc3_0, 
							fps_tpl_irq_ttc2_2, 
							fps_tpl_irq_ttc2_1, 
							fps_tpl_irq_ttc2_0, 
							fps_tpl_irq_ttc1_2, 
							fps_tpl_irq_ttc1_1, 
							fps_tpl_irq_ttc1_0, 
							fps_tpl_irq_ttc0_2, 
							fps_tpl_irq_ttc0_1, 
							fps_tpl_irq_ttc0_0, 
							fps_tpl_irq_ipi_channel0, 
							fps_tpl_irq_ipi_channel1, 
							fps_tpl_irq_ipi_channel2, 
							fps_tpl_irq_ipi_channel7, 
							fps_tpl_irq_ipi_channel8, 
							fps_tpl_irq_ipi_channel9, 
							fps_tpl_irq_ipi_channel10, 
							fps_tpl_irq_clkmon, 
							fps_tpl_irq_rtc_seconds, 
							fps_tpl_irq_rtc_alaram, 
							fps_tpl_irq_lpd_apm, 
							fps_tpl_irq_can1, 
							fps_tpl_irq_can0, 
							fps_tpl_irq_uart1, 
							fps_tpl_irq_uart0, 
							fps_tpl_irq_spi1, 
							fps_tpl_irq_spi0, 
							fps_tpl_irq_i2c1, 
							fps_tpl_irq_i2c0, 
							fps_tpl_irq_gpio, 
							fps_tpl_irq_qspi, 
							fps_tpl_irq_nand, 
							fps_tpl_irq_r5_core1_ecc_error, 
							fps_tpl_irq_r5_core0_ecc_error, 
							fps_tpl_irq_lpd_apb_intr, 
							fps_tpl_irq_ocm_error, 
							fps_tpl_irq_rpu_pm, 
							irq_lpd_dev_null[7:0]}),
.PSPLIRQFPD ({irq_fpd_dev_null[19:12], 
							fps_tpl_irq_intf_fpd_smmu, 
							fps_tpl_irq_intf_ppd_cci, 
							fps_tpl_irq_apu_regs, 
							fps_tpl_irq_apu_exterr, 
							fps_tpl_irq_apu_l2err, 
							fps_tpl_irq_apu_comm, 
							fps_tpl_irq_apu_pmu, 
							fps_tpl_irq_apu_cti, 
							fps_tpl_irq_apu_cpumnt, 
							fps_tpl_irq_xmpu_fpd, 
							fps_tpl_irq_sata, 
							fps_tpl_irq_gpu, 
							fps_tpl_irq_gdma_chan, 
							fps_tpl_irq_apm_fpd, 
							fps_tpl_irq_dpdma, 
							fps_tpl_irq_fpd_atb_error, 
							fps_tpl_irq_fpd_apb_int, 
							fps_tpl_irq_dport, 
							fps_tpl_irq_pcie_msc, 
							fps_tpl_irq_pcie_dma, 
							fps_tpl_irq_pcie_legacy, 
							fps_tpl_irq_pcie_msi, 
							fps_tpl_irq_fp_wdt, 
							fps_tpl_irq_ddr_ss, 
							irq_fpd_dev_null[11:0]}),
.OSCRTCCLK (osc_rtc_clk),
.PLPMUGPI (pl_pmu_gpi),
.PMUPLGPO (pmu_pl_gpo),
.AIBPMUAFIFMFPDACK (aib_pmu_afifm_fpd_ack),
.AIBPMUAFIFMLPDACK (aib_pmu_afifm_lpd_ack),
.PMUAIBAFIFMFPDREQ (pmu_aib_afifm_fpd_req),
.PMUAIBAFIFMLPDREQ (pmu_aib_afifm_lpd_req),
.PMUERRORTOPL (pmu_error_to_pl),
.PMUERRORFROMPL (pmu_error_from_pl),
.DDRCEXTREFRESHRANK0REQ (ddrc_ext_refresh_rank0_req),
.DDRCEXTREFRESHRANK1REQ (ddrc_ext_refresh_rank1_req),
.DDRCREFRESHPLCLK (clk_tps_fpl_ddrc_refresh),
.PLACPINACT (pl_acpinact),
.PLCLK (clk_fps_tpl_clks),
.DPVIDEOREFCLK(clk_fps_tpl_dp_video),
.DPAUDIOREFCLK(clk_fps_tpl_dp_audio),
.PSS_ALTO_CORE_PAD_MGTTXN0OUT(pss_alto_core_pad_mgttxn0out),// What are these?
.PSS_ALTO_CORE_PAD_MGTTXN1OUT(pss_alto_core_pad_mgttxn1out),
.PSS_ALTO_CORE_PAD_MGTTXN2OUT(pss_alto_core_pad_mgttxn2out),
.PSS_ALTO_CORE_PAD_MGTTXN3OUT(pss_alto_core_pad_mgttxn3out),
.PSS_ALTO_CORE_PAD_MGTTXP0OUT(pss_alto_core_pad_mgttxp0out),
.PSS_ALTO_CORE_PAD_MGTTXP1OUT(pss_alto_core_pad_mgttxp1out),
.PSS_ALTO_CORE_PAD_MGTTXP2OUT(pss_alto_core_pad_mgttxp2out),
.PSS_ALTO_CORE_PAD_MGTTXP3OUT(pss_alto_core_pad_mgttxp3out),
.PSS_ALTO_CORE_PAD_PADO(pss_alto_core_pad_pad0),
.PSS_ALTO_CORE_PAD_BOOTMODE(),
.PSS_ALTO_CORE_PAD_CLK(),
.PSS_ALTO_CORE_PAD_DONEB(),
.PSS_ALTO_CORE_PAD_DRAMA(),
.PSS_ALTO_CORE_PAD_DRAMACTN(),
.PSS_ALTO_CORE_PAD_DRAMALERTN(),
.PSS_ALTO_CORE_PAD_DRAMBA(),
.PSS_ALTO_CORE_PAD_DRAMBG(),
.PSS_ALTO_CORE_PAD_DRAMCK(),
.PSS_ALTO_CORE_PAD_DRAMCKE(),
.PSS_ALTO_CORE_PAD_DRAMCKN(),
.PSS_ALTO_CORE_PAD_DRAMCSN(),
.PSS_ALTO_CORE_PAD_DRAMDM(),
.PSS_ALTO_CORE_PAD_DRAMDQ(),
.PSS_ALTO_CORE_PAD_DRAMDQS(),
.PSS_ALTO_CORE_PAD_DRAMDQSN(),
.PSS_ALTO_CORE_PAD_DRAMODT(),
.PSS_ALTO_CORE_PAD_DRAMPARITY(),
.PSS_ALTO_CORE_PAD_DRAMRAMRSTN(),
.PSS_ALTO_CORE_PAD_ERROROUT(),
.PSS_ALTO_CORE_PAD_ERRORSTATUS(),
.PSS_ALTO_CORE_PAD_INITB(),
.PSS_ALTO_CORE_PAD_JTAGTCK(),
.PSS_ALTO_CORE_PAD_JTAGTDI(),
.PSS_ALTO_CORE_PAD_JTAGTDO(),
.PSS_ALTO_CORE_PAD_JTAGTMS(),
.PSS_ALTO_CORE_PAD_MIO(),
.PSS_ALTO_CORE_PAD_PORB(),
.PSS_ALTO_CORE_PAD_PROGB(),
.PSS_ALTO_CORE_PAD_RCALIBINOUT(),
.PSS_ALTO_CORE_PAD_SRSTB(),
.PSS_ALTO_CORE_PAD_ZQ(),
.PSS_ALTO_CORE_PAD_MGTRXN0IN(),
.PSS_ALTO_CORE_PAD_MGTRXN1IN(),
.PSS_ALTO_CORE_PAD_MGTRXN2IN(),
.PSS_ALTO_CORE_PAD_MGTRXN3IN(),
.PSS_ALTO_CORE_PAD_MGTRXP0IN(),
.PSS_ALTO_CORE_PAD_MGTRXP1IN(),
.PSS_ALTO_CORE_PAD_MGTRXP2IN(),
.PSS_ALTO_CORE_PAD_MGTRXP3IN(),
.PSS_ALTO_CORE_PAD_PADI(),
.PSS_ALTO_CORE_PAD_REFN0IN(),
.PSS_ALTO_CORE_PAD_REFN1IN(),
.PSS_ALTO_CORE_PAD_REFN2IN(),
.PSS_ALTO_CORE_PAD_REFN3IN(),
.PSS_ALTO_CORE_PAD_REFP0IN(),
.PSS_ALTO_CORE_PAD_REFP1IN(),
.PSS_ALTO_CORE_PAD_REFP2IN(),
.PSS_ALTO_CORE_PAD_REFP3IN()
);

endmodule

